--------------------------------------------------------------------------------
--                         ModuloCounter_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_28_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of ModuloCounter_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(4 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 27 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1356461_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1356463)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1356461_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1356461_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1356466
--                  (IntAdderAlternative_27_f250_uid1356470)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1356466 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1356466 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1356473
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1356473 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1356473 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1356476
--                   (IntAdderClassical_34_f250_uid1356478)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1356476 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1356476 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1356461
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1356461 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1356461 is
   component FPAdd_8_23_uid1356461_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1356466 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1356473 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1356476 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1356461_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1356466  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1356473  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1356476  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1356461 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1356461  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_28_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
         iS_23 when "10111",
         iS_24 when "11000",
         iS_25 when "11001",
         iS_26 when "11010",
         iS_27 when "11011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1357122
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1357122 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1357122 is
signal XX_m1357123 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1357123 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1357123 <= X ;
   YY_m1357123 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1357126
--                   (IntAdderClassical_33_f500_uid1357128)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1357126 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1357126 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1357122 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1357126 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1357122  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid1357126  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1357385_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1357387)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1357385_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1357385_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1357390
--                  (IntAdderAlternative_27_f250_uid1357394)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1357390 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1357390 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1357397
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1357397 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1357397 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1357400
--                   (IntAdderClassical_34_f250_uid1357402)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1357400 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1357400 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1357385
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1357385 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1357385 is
   component FPAdd_8_23_uid1357385_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1357390 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1357397 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1357400 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1357385_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1357390  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1357397  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1357400  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid1357385 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid1357385  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_23_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_23_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "001" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "010" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "011" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "100" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "001" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "010" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "011" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "100" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "011" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "100" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "001" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "010" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "011" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "100" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "001" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "010" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "001" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "010" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "011" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "100" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "001" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "010" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "011" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "100" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "011" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "100" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "001" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "010" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "010" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "011" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "100" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "001" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "010" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "011" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "100" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "001" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "001" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "010" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "011" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "100" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "001" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "010" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "011" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "100" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "011" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "100" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "001" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "010" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "011" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "100" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "001" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "010" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "001" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "010" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "011" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "100" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "001" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "010" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "011" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "100" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "011" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "100" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "001" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "010" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "001" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "010" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "011" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "100" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "001" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "010" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "011" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "100" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "011" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "100" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "001" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "010" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "011" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "100" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "001" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "010" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "001" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "010" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "011" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "100" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "010" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "011" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "100" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "001" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "011" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "100" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "001" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "010" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "001" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "010" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "011" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "100" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "001" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "010" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "011" when "10101",
      "000" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "100" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "000" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "011" when "00101",
      "000" when "00110",
      "000" when "00111",
      "000" when "01000",
      "000" when "01001",
      "100" when "01010",
      "000" when "01011",
      "000" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "001" when "10110",
      "000" when "10111",
      "000" when "11000",
      "000" when "11001",
      "000" when "11010",
      "010" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "000" when "00000",
      "010" when "00001",
      "000" when "00010",
      "000" when "00011",
      "000" when "00100",
      "000" when "00101",
      "000" when "00110",
      "011" when "00111",
      "000" when "01000",
      "000" when "01001",
      "000" when "01010",
      "000" when "01011",
      "100" when "01100",
      "000" when "01101",
      "000" when "01110",
      "000" when "01111",
      "000" when "10000",
      "000" when "10001",
      "000" when "10010",
      "000" when "10011",
      "000" when "10100",
      "000" when "10101",
      "000" when "10110",
      "000" when "10111",
      "001" when "11000",
      "000" when "11001",
      "000" when "11010",
      "000" when "11011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "01010" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "01000" when "00011",
      "01001" when "00100",
      "01011" when "00101",
      "00000" when "00110",
      "00111" when "00111",
      "10110" when "01000",
      "00101" when "01001",
      "00110" when "01010",
      "10010" when "01011",
      "00000" when "01100",
      "10001" when "01101",
      "10100" when "01110",
      "10101" when "01111",
      "00100" when "10000",
      "00000" when "10001",
      "00010" when "10010",
      "10011" when "10011",
      "00011" when "10100",
      "00001" when "10101",
      "01110" when "10110",
      "00000" when "10111",
      "01101" when "11000",
      "01100" when "11001",
      "01111" when "11010",
      "10000" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "01110" when "00000",
      "00000" when "00001",
      "01010" when "00010",
      "10110" when "00011",
      "01101" when "00100",
      "01001" when "00101",
      "00000" when "00110",
      "10010" when "00111",
      "00100" when "01000",
      "10100" when "01001",
      "10101" when "01010",
      "00111" when "01011",
      "00000" when "01100",
      "00010" when "01101",
      "00011" when "01110",
      "01000" when "01111",
      "10011" when "10000",
      "00000" when "10001",
      "01111" when "10010",
      "00110" when "10011",
      "10000" when "10100",
      "10001" when "10101",
      "01100" when "10110",
      "00000" when "10111",
      "01011" when "11000",
      "00000" when "11001",
      "00101" when "11010",
      "00001" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "10110" when "00000",
      "00000" when "00001",
      "00001" when "00010",
      "10101" when "00011",
      "10000" when "00100",
      "01000" when "00101",
      "00000" when "00110",
      "01111" when "00111",
      "10100" when "01000",
      "10001" when "01001",
      "10011" when "01010",
      "01100" when "01011",
      "00000" when "01100",
      "01011" when "01101",
      "00000" when "01110",
      "10010" when "01111",
      "01101" when "10000",
      "00000" when "10001",
      "00011" when "10010",
      "01110" when "10011",
      "00111" when "10100",
      "00010" when "10101",
      "00110" when "10110",
      "00000" when "10111",
      "00101" when "11000",
      "00100" when "11001",
      "01001" when "11010",
      "01010" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00111" when "00000",
      "00000" when "00001",
      "01011" when "00010",
      "00110" when "00011",
      "00100" when "00100",
      "00010" when "00101",
      "00000" when "00110",
      "00011" when "00111",
      "00101" when "01000",
      "10010" when "01001",
      "10011" when "01010",
      "10000" when "01011",
      "00000" when "01100",
      "01101" when "01101",
      "10110" when "01110",
      "10001" when "01111",
      "01111" when "10000",
      "00000" when "10001",
      "01010" when "10010",
      "01110" when "10011",
      "01100" when "10100",
      "01001" when "10101",
      "10101" when "10110",
      "00000" when "10111",
      "10100" when "11000",
      "00000" when "11001",
      "01000" when "11010",
      "00001" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00010" when "00000",
      "00000" when "00001",
      "00101" when "00010",
      "00001" when "00011",
      "00000" when "00100",
      "01010" when "00101",
      "00000" when "00110",
      "01110" when "00111",
      "10110" when "01000",
      "10001" when "01001",
      "10011" when "01010",
      "10000" when "01011",
      "00000" when "01100",
      "01101" when "01101",
      "10010" when "01110",
      "10101" when "01111",
      "10100" when "10000",
      "00000" when "10001",
      "00110" when "10010",
      "01111" when "10011",
      "01001" when "10100",
      "00011" when "10101",
      "01000" when "10110",
      "00000" when "10111",
      "00111" when "11000",
      "00100" when "11001",
      "01011" when "11010",
      "01100" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "10110" when "00000",
      "00000" when "00001",
      "00001" when "00010",
      "10101" when "00011",
      "10100" when "00100",
      "00010" when "00101",
      "00000" when "00110",
      "00011" when "00111",
      "00101" when "01000",
      "01100" when "01001",
      "10000" when "01010",
      "01101" when "01011",
      "00000" when "01100",
      "01010" when "01101",
      "01011" when "01110",
      "01111" when "01111",
      "01110" when "10000",
      "00000" when "10001",
      "00111" when "10010",
      "01001" when "10011",
      "01000" when "10100",
      "10011" when "10101",
      "10010" when "10110",
      "00000" when "10111",
      "10001" when "11000",
      "00110" when "11001",
      "00100" when "11010",
      "00000" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "10101" when "00000",
      "00000" when "00001",
      "00010" when "00010",
      "10100" when "00011",
      "10011" when "00100",
      "10010" when "00101",
      "00000" when "00110",
      "10001" when "00111",
      "10110" when "01000",
      "00110" when "01001",
      "01000" when "01010",
      "01111" when "01011",
      "00000" when "01100",
      "01101" when "01101",
      "00101" when "01110",
      "00111" when "01111",
      "10000" when "10000",
      "00000" when "10001",
      "00011" when "10010",
      "01110" when "10011",
      "00100" when "10100",
      "01100" when "10101",
      "01010" when "10110",
      "00000" when "10111",
      "01001" when "11000",
      "01011" when "11001",
      "00001" when "11010",
      "00000" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00101" when "00000",
      "00000" when "00001",
      "10110" when "00010",
      "00011" when "00011",
      "00010" when "00100",
      "00001" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00100" when "01000",
      "10010" when "01001",
      "10100" when "01010",
      "01011" when "01011",
      "00000" when "01100",
      "01001" when "01101",
      "10011" when "01110",
      "10101" when "01111",
      "01010" when "10000",
      "00000" when "10001",
      "01100" when "10010",
      "01000" when "10011",
      "01111" when "10100",
      "00111" when "10101",
      "01110" when "10110",
      "00000" when "10111",
      "01101" when "11000",
      "00110" when "11001",
      "10000" when "11010",
      "10001" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_28_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(4 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_28_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_23_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount281_out : std_logic_vector(4 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product316_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product316_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product213_4_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product213_4_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product316_4_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product316_4_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No20_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No21_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No22_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No23_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No3_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No24_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No10_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No11_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No12_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No13_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No14_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Subtract16_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Subtract16_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No25_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Subtract16_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Subtract16_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No26_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No1_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Subtract16_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Subtract16_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No2_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Subtract16_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Subtract16_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No28_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No3_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Subtract16_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Subtract16_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No29_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No4_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product316_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product316_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product316_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product316_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No1_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No1_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No2_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No2_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No3_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No4_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay74No4_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount281_instance: ModuloCounter_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount281_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg32_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg40_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg56_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg56_out;
SharedReg64_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg48_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg72_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg83_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
SharedReg94_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg105_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg116_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg127_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg151_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg163_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg175_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg187_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg205_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg223_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg223_out;
SharedReg241_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg259_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg223_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg32_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg40_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg56_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg56_out;
SharedReg64_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg72_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
SharedReg94_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg105_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg116_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg187_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg205_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg223_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg223_out;
SharedReg241_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg259_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg223_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg151_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg72_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg83_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
SharedReg94_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg105_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg116_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg40_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg48_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg56_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg56_out;
SharedReg64_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg64_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg48_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg72_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg83_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
SharedReg94_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg116_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg127_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg151_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg175_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg139_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg151_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg163_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg175_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg205_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg223_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg223_out;
SharedReg241_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg259_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg223_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg187_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg205_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg223_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg223_out;
SharedReg241_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg259_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg223_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg127_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg139_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg151_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg163_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg175_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg163_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg699_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg709_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg719_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg729_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg719_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg803_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg767_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg791_out;
SharedReg815_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg767_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg779_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg791_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg767_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg567_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg581_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg581_out;
SharedReg595_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg595_out;
SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg609_out;
SharedReg623_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg623_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg581_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg595_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg623_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg372_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg388_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg404_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg420_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg436_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg436_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg436_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg372_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg388_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg404_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg420_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg436_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg436_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg436_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg699_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg709_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg719_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg729_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg719_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg767_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg767_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg699_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg709_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg719_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg729_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg719_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg699_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg709_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg719_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg729_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg719_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg767_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg581_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg581_out;
SharedReg595_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg595_out;
SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg609_out;
SharedReg623_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg623_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg581_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg595_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg623_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg699_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg709_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg719_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg729_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg719_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg767_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg767_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg779_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg791_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg803_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg803_out;
SharedReg815_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg791_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg803_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg573_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg278_out;
SharedReg575_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg575_out;
SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg136_out;
SharedReg386_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg386_out;
SharedReg384_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg384_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg567_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg769_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg769_out;
SharedReg375_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg375_out;
SharedReg316_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg316_out;
SharedReg196_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg196_out;
SharedReg131_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg131_out;
SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg278_out;
SharedReg458_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg458_out;
SharedReg767_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg767_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg567_out;
SharedReg373_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg373_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg567_out;
SharedReg699_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg699_out;
SharedReg318_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg318_out;
SharedReg133_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg133_out;
SharedReg381_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg381_out;
SharedReg195_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg195_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg769_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg375_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg316_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg196_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg131_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg458_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg767_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg373_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg699_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg318_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg133_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg381_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg195_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg278_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg575_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg136_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg386_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg384_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg578_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg578_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg317_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg317_out;
SharedReg377_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg377_out;
SharedReg75_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg75_out;
SharedReg378_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg378_out;
SharedReg573_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg573_out;
SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg699_out;
SharedReg767_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg767_out;
SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg699_out;
SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
SharedReg452_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg452_out;
SharedReg204_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg204_out;
SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg187_out;
SharedReg316_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg316_out;
SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg277_out;
SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg372_out;
SharedReg383_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg383_out;
SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg372_out;
SharedReg769_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg769_out;
SharedReg373_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg373_out;
SharedReg505_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg505_out;
SharedReg74_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg74_out;
SharedReg570_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg570_out;
SharedReg130_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg130_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg578_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg767_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg699_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg452_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg204_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg316_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg383_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg372_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg769_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg373_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg505_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg74_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg570_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg130_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg317_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg377_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg75_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg378_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg573_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg709_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg328_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg328_out;
SharedReg145_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg397_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg397_out;
SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg213_out;
SharedReg587_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg587_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg284_out;
SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg589_out;
SharedReg148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg148_out;
SharedReg402_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg402_out;
SharedReg400_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg400_out;
SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg581_out;
SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg581_out;
SharedReg781_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg781_out;
SharedReg391_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg391_out;
SharedReg326_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg326_out;
SharedReg214_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg214_out;
SharedReg143_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg143_out;
SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg284_out;
SharedReg468_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg468_out;
SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg779_out;
SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg581_out;
SharedReg389_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg389_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg402_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg400_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg781_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg391_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg328_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg326_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg214_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg143_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg284_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg468_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg389_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg145_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg397_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg587_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg781_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg781_out;
SharedReg389_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg514_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg514_out;
SharedReg85_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg85_out;
SharedReg584_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg584_out;
SharedReg142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg142_out;
SharedReg592_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg592_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg327_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg327_out;
SharedReg393_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg393_out;
SharedReg86_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg86_out;
SharedReg394_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg394_out;
SharedReg587_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg587_out;
SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg709_out;
SharedReg779_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg779_out;
SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg709_out;
SharedReg582_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg582_out;
SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg462_out;
SharedReg222_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg222_out;
SharedReg205_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg205_out;
SharedReg326_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg326_out;
SharedReg283_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg283_out;
SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg388_out;
SharedReg399_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg399_out;
SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg388_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg781_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg327_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg393_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg86_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg394_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg587_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg779_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg709_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg582_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg514_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg222_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg205_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg326_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg283_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg399_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg388_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg85_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg584_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg592_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg514_out;
SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg478_out;
SharedReg791_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg595_out;
SharedReg405_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg405_out;
SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg719_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg719_out;
SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg547_out;
SharedReg157_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg157_out;
SharedReg413_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg413_out;
SharedReg231_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg231_out;
SharedReg601_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg601_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg2_out;
SharedReg290_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg290_out;
SharedReg603_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg603_out;
SharedReg160_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg160_out;
SharedReg418_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg418_out;
SharedReg416_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg416_out;
SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg595_out;
SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg595_out;
SharedReg793_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg793_out;
SharedReg407_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg407_out;
SharedReg336_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg336_out;
SharedReg232_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg232_out;
SharedReg155_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg155_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg231_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg601_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg290_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg603_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg160_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg418_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg791_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg416_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg793_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg407_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg336_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg232_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg155_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg405_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg719_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg157_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg413_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg336_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg289_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg289_out;
SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg415_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg415_out;
SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg404_out;
SharedReg793_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg793_out;
SharedReg405_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
SharedReg296_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg296_out;
SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg96_out;
SharedReg598_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg598_out;
SharedReg154_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg154_out;
SharedReg606_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg606_out;
SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg18_out;
SharedReg337_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg337_out;
SharedReg409_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg409_out;
SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg97_out;
SharedReg410_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg410_out;
SharedReg601_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg601_out;
SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg719_out;
SharedReg791_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg791_out;
SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg719_out;
SharedReg596_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg596_out;
SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg472_out;
SharedReg240_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg240_out;
SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg223_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg289_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg154_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg606_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg337_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg409_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg410_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg601_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg791_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg719_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg596_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg240_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg415_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg404_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg793_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg296_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg598_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg805_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg805_out;
SharedReg423_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg423_out;
SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg362_out;
SharedReg250_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg250_out;
SharedReg167_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg167_out;
SharedReg296_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg296_out;
SharedReg488_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg488_out;
SharedReg803_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg803_out;
SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg609_out;
SharedReg421_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg421_out;
SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg609_out;
SharedReg729_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg729_out;
SharedReg364_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg364_out;
SharedReg169_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg169_out;
SharedReg429_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg429_out;
SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg249_out;
SharedReg615_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg615_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg2_out;
SharedReg311_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg311_out;
SharedReg617_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg617_out;
SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg172_out;
SharedReg434_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg434_out;
SharedReg432_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg432_out;
SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg609_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg805_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg421_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg729_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg364_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg169_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg429_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg615_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg423_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg311_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg617_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg434_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg432_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg250_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg167_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg296_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg488_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg803_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg609_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg803_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg729_out;
SharedReg610_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg610_out;
SharedReg482_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg482_out;
SharedReg258_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg258_out;
SharedReg241_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg241_out;
SharedReg362_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg362_out;
SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg310_out;
SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg420_out;
SharedReg431_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg431_out;
SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg420_out;
SharedReg805_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg805_out;
SharedReg421_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg421_out;
SharedReg523_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg523_out;
SharedReg107_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg107_out;
SharedReg612_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg612_out;
SharedReg166_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg166_out;
SharedReg620_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg620_out;
SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg18_out;
SharedReg363_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg363_out;
SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg425_out;
SharedReg108_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg108_out;
SharedReg426_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg426_out;
SharedReg615_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg615_out;
SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg729_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg805_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg421_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg523_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg107_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg612_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg166_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg620_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg610_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg363_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg108_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg426_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg615_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg729_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg482_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg258_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg241_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg362_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg420_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg431_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg631_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg631_out;
SharedReg184_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg184_out;
SharedReg450_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg450_out;
SharedReg448_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg448_out;
SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg623_out;
SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg623_out;
SharedReg817_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg817_out;
SharedReg439_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg439_out;
SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg353_out;
SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg268_out;
SharedReg179_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg179_out;
SharedReg523_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg523_out;
SharedReg499_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg499_out;
SharedReg815_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg815_out;
SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg623_out;
SharedReg437_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg437_out;
SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg623_out;
SharedReg739_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg739_out;
SharedReg554_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg554_out;
SharedReg181_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg181_out;
SharedReg445_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg445_out;
SharedReg267_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg267_out;
SharedReg629_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg629_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg2_out;
SharedReg305_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg305_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg631_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg179_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg523_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg499_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg815_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg437_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg739_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg554_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg181_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg450_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg445_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg267_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg629_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg305_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg448_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg623_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg817_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg439_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg441_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg441_out;
SharedReg119_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg119_out;
SharedReg442_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg442_out;
SharedReg629_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg629_out;
SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg739_out;
SharedReg815_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg815_out;
SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg739_out;
SharedReg624_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg624_out;
SharedReg493_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg493_out;
SharedReg276_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg276_out;
SharedReg259_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg259_out;
SharedReg353_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg353_out;
SharedReg304_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg304_out;
SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg436_out;
SharedReg447_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg447_out;
SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg436_out;
SharedReg817_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg817_out;
SharedReg437_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg437_out;
SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg531_out;
SharedReg118_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg118_out;
SharedReg626_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg626_out;
SharedReg178_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg178_out;
SharedReg634_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg634_out;
SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg18_out;
SharedReg354_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg354_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg441_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg259_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg353_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg304_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg447_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg436_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg817_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg437_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg118_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg442_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg626_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg178_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg634_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg354_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg629_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg815_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg739_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg624_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg493_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg276_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg452_out;
SharedReg316_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg316_out;
SharedReg277_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg277_out;
SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg198_out;
SharedReg572_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg572_out;
SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg72_out;
SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg72_out;
SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg189_out;
SharedReg35_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg35_out;
SharedReg321_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg321_out;
SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg452_out;
SharedReg776_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg776_out;
SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg452_out;
SharedReg323_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg323_out;
SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg188_out;
SharedReg128_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg73_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg73_out;
SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg72_out;
SharedReg187_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg187_out;
SharedReg506_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg506_out;
Delay19No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast <= Delay19No_out;
SharedReg687_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg687_out;
SharedReg382_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg382_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg189_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg35_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg321_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg776_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg323_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg188_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg73_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg72_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg187_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg506_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay19No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg687_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg382_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg10_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg452_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg316_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg277_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg572_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No42_out);

SharedReg39_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg504_out;
SharedReg750_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg750_out;
SharedReg320_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg320_out;
SharedReg132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg132_out;
SharedReg580_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg580_out;
SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg187_out;
SharedReg128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg128_out;
SharedReg282_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg282_out;
SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg504_out;
SharedReg778_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg778_out;
SharedReg687_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg687_out;
SharedReg316_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg316_out;
SharedReg32_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg32_out;
SharedReg82_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg82_out;
SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg127_out;
SharedReg188_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg188_out;
SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg33_out;
SharedReg319_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg319_out;
SharedReg318_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg318_out;
SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg539_out;
SharedReg574_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg574_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg282_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg778_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg687_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg316_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg32_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg82_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg127_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg188_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg319_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg318_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg574_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg504_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg750_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg320_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg580_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg515_out;
Delay19No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= Delay19No1_out;
SharedReg647_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg647_out;
SharedReg398_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg398_out;
SharedReg146_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg146_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg462_out;
SharedReg326_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg326_out;
SharedReg283_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg283_out;
SharedReg216_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg216_out;
SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg586_out;
SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg83_out;
SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg83_out;
SharedReg207_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg207_out;
SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg43_out;
SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg331_out;
SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg462_out;
SharedReg788_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg788_out;
SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg462_out;
SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg333_out;
SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg206_out;
SharedReg140_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg140_out;
SharedReg84_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg84_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg326_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg283_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg216_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg83_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg207_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg788_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg462_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg140_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg84_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay19No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg647_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg398_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg146_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg10_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No44_out);

SharedReg206_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg41_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg541_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg541_out;
SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg546_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg546_out;
SharedReg588_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg588_out;
SharedReg47_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg47_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg513_out;
SharedReg660_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg660_out;
SharedReg330_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg330_out;
SharedReg144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg144_out;
SharedReg594_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg594_out;
SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg139_out;
SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg205_out;
SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg205_out;
SharedReg140_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg140_out;
SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg288_out;
SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg513_out;
SharedReg790_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg790_out;
SharedReg647_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg647_out;
SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg326_out;
SharedReg40_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg40_out;
SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg93_out;
SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg139_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg660_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg330_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg594_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg140_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg541_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg513_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg790_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg647_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg40_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg546_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg588_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg47_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg472_out;
SharedReg343_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg343_out;
SharedReg224_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg224_out;
SharedReg152_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg223_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg223_out;
SharedReg661_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg661_out;
Delay19No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= Delay19No2_out;
SharedReg654_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg654_out;
SharedReg414_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg414_out;
SharedReg158_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg158_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg12_out;
SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg472_out;
SharedReg336_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg336_out;
SharedReg289_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg289_out;
SharedReg234_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg234_out;
SharedReg600_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg600_out;
SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg94_out;
SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg94_out;
SharedReg225_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg225_out;
SharedReg51_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg51_out;
SharedReg341_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg341_out;
SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg472_out;
SharedReg800_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg800_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg343_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg414_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg158_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg336_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg289_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg234_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg224_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg600_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg225_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg51_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg341_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg472_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg800_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg152_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg223_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg661_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay19No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg654_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No46_out);

SharedReg654_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg654_out;
SharedReg336_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg336_out;
SharedReg48_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg104_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg104_out;
SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg151_out;
SharedReg224_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg224_out;
SharedReg49_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg49_out;
SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg339_out;
SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg338_out;
SharedReg347_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg347_out;
SharedReg602_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg602_out;
SharedReg55_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg55_out;
SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg28_out;
SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg295_out;
SharedReg669_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg669_out;
SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg340_out;
SharedReg156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg156_out;
SharedReg608_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg608_out;
SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg151_out;
SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg223_out;
SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg223_out;
SharedReg152_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg152_out;
SharedReg294_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg294_out;
SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg295_out;
SharedReg802_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg802_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg654_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg602_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg55_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg669_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg48_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg608_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg152_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg294_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg295_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg802_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg104_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg151_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg224_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg49_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg347_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg243_out;
SharedReg59_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg367_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg367_out;
SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg482_out;
SharedReg812_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg812_out;
SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg482_out;
SharedReg369_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg369_out;
SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg242_out;
SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg164_out;
SharedReg106_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg106_out;
SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg105_out;
SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg241_out;
SharedReg524_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg524_out;
Delay19No3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast <= Delay19No3_out;
SharedReg639_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg639_out;
SharedReg430_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg430_out;
SharedReg170_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg170_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg12_out;
SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg482_out;
SharedReg362_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg362_out;
SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg310_out;
SharedReg252_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg252_out;
SharedReg614_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg614_out;
SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg105_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg106_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg524_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay19No3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg639_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg430_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg170_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg59_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg362_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg252_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg614_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg105_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg367_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg812_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg369_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No48_out);

SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg241_out;
SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg241_out;
SharedReg164_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg164_out;
SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg315_out;
SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg522_out;
SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg814_out;
SharedReg639_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg639_out;
SharedReg362_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg56_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg56_out;
SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg115_out;
SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg163_out;
SharedReg242_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg242_out;
SharedReg57_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg57_out;
SharedReg349_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg349_out;
SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg364_out;
SharedReg553_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg553_out;
SharedReg616_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg616_out;
SharedReg63_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg63_out;
SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg28_out;
SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg522_out;
SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg678_out;
SharedReg366_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg366_out;
SharedReg168_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg168_out;
SharedReg622_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg622_out;
SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg163_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg242_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg57_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg349_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg553_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg616_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg63_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg164_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg366_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg168_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg622_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg163_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg522_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg639_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg56_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg304_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg304_out;
SharedReg270_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg270_out;
SharedReg628_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg628_out;
SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg261_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg67_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg67_out;
SharedReg358_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg358_out;
SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg493_out;
SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg824_out;
SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg493_out;
SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg260_out;
SharedReg176_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg176_out;
SharedReg117_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg117_out;
SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg116_out;
SharedReg259_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg259_out;
SharedReg679_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg679_out;
Delay19No4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast <= Delay19No4_out;
SharedReg694_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg694_out;
SharedReg446_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg446_out;
SharedReg182_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg182_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg12_out;
SharedReg637_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg637_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg304_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg176_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg259_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg679_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay19No4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg270_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg694_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg446_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg182_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg637_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg628_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg67_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg358_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg493_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No50_out);

SharedReg494_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg494_out;
SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg180_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg180_out;
SharedReg636_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg259_out;
SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg259_out;
SharedReg176_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg176_out;
SharedReg309_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg309_out;
SharedReg530_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg530_out;
SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg826_out;
SharedReg694_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg694_out;
SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg353_out;
SharedReg64_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg64_out;
SharedReg126_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg126_out;
SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg175_out;
SharedReg260_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg260_out;
SharedReg65_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg65_out;
SharedReg356_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg356_out;
SharedReg355_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg355_out;
SharedReg561_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg561_out;
SharedReg630_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg630_out;
SharedReg71_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg71_out;
SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg28_out;
SharedReg677_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg677_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg494_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg64_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg126_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg260_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg65_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg356_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg355_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg180_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg561_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg630_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg71_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg677_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg636_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg259_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg176_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg309_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg530_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No52_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg316_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg7_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg319_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg319_out;
SharedReg538_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg538_out;
SharedReg456_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg456_out;
SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg377_out;
SharedReg76_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg76_out;
SharedReg133_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg133_out;
SharedReg194_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg194_out;
SharedReg277_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg277_out;
SharedReg279_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg279_out;
SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg460_out;
SharedReg543_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg543_out;
SharedReg458_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg458_out;
SharedReg541_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg541_out;
SharedReg755_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg755_out;
SharedReg706_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg706_out;
SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg316_out;
SharedReg700_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg700_out;
SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg377_out;
SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg377_out;
SharedReg540_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg540_out;
SharedReg691_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg691_out;
SharedReg278_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg278_out;
SharedReg80_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg80_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg133_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg194_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg277_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg279_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg543_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg458_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg541_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg755_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg706_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg6_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg316_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg700_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg540_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg691_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg278_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg80_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg319_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg538_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg456_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg76_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No52_out);

SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg452_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg23_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg455_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg455_out;
SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg685_out;
SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg538_out;
SharedReg387_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg387_out;
SharedReg199_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg199_out;
SharedReg138_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg138_out;
SharedReg202_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg202_out;
SharedReg318_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg318_out;
SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg316_out;
SharedReg459_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg459_out;
SharedReg690_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg690_out;
SharedReg504_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg504_out;
SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg685_out;
SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg538_out;
SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg699_out;
SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg452_out;
SharedReg708_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg708_out;
SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg699_out;
SharedReg372_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg372_out;
SharedReg541_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg541_out;
SharedReg317_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg317_out;
SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg316_out;
SharedReg78_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg78_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg138_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg318_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg459_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg690_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg504_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg22_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg452_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg708_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg699_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg372_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg541_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg317_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg316_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg78_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg455_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg685_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg538_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg387_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg199_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No54_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg393_out;
SharedReg547_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg651_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg651_out;
SharedReg284_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg91_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg91_out;
SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg326_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg7_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg329_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg329_out;
SharedReg545_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg545_out;
SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg466_out;
SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg393_out;
SharedReg87_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg87_out;
SharedReg145_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg145_out;
SharedReg212_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg212_out;
SharedReg283_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg283_out;
SharedReg285_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg285_out;
SharedReg470_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg470_out;
SharedReg550_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg550_out;
SharedReg468_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg468_out;
SharedReg548_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg548_out;
SharedReg665_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg665_out;
SharedReg716_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg716_out;
SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg326_out;
SharedReg710_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg710_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg329_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg545_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg393_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg87_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg145_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg212_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg283_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg285_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg547_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg470_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg550_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg468_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg548_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg665_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg716_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg710_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg651_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg91_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No54_out);

SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg709_out;
SharedReg388_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg286_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg327_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg327_out;
SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg89_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg462_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg23_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg465_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg465_out;
SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg645_out;
SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg545_out;
SharedReg403_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg403_out;
SharedReg217_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg217_out;
SharedReg150_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg150_out;
SharedReg220_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg220_out;
SharedReg328_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg328_out;
SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg326_out;
SharedReg469_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg469_out;
SharedReg650_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg650_out;
SharedReg513_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg513_out;
SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg645_out;
SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg545_out;
SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg709_out;
SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg462_out;
SharedReg718_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg718_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg465_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg403_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg217_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg150_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg220_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg328_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg286_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg469_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg650_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg513_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg645_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg545_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg709_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg718_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg327_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg462_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_2_impl_out,
                 X => Delay1No56_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg349_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg674_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg674_out;
SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg726_out;
SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg336_out;
SharedReg720_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg720_out;
SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg409_out;
SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg291_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg658_out;
SharedReg290_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg290_out;
SharedReg102_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg102_out;
SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg336_out;
SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg11_out;
SharedReg7_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg7_out;
SharedReg339_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg339_out;
SharedReg346_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg346_out;
SharedReg476_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg476_out;
SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg409_out;
SharedReg98_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg98_out;
SharedReg157_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg157_out;
SharedReg230_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg230_out;
SharedReg289_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg289_out;
SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg291_out;
SharedReg480_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg480_out;
SharedReg351_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg351_out;
SharedReg478_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg478_out;
   MUX_Add12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg674_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg102_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg7_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg339_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg346_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg476_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg98_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg157_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg230_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg289_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg480_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg351_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg478_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg336_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg720_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg409_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg291_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg290_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_2_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_0_out,
                 Y => Delay1No56_out);

SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg472_out;
SharedReg728_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg728_out;
SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg719_out;
SharedReg404_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg404_out;
SharedReg349_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg349_out;
SharedReg337_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg337_out;
SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg336_out;
SharedReg100_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg100_out;
SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg472_out;
SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg23_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg23_out;
SharedReg475_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg475_out;
SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg652_out;
SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg346_out;
SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg419_out;
SharedReg235_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg235_out;
SharedReg162_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg162_out;
SharedReg238_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg238_out;
SharedReg338_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg338_out;
SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg336_out;
SharedReg479_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg479_out;
SharedReg657_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg657_out;
SharedReg659_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg659_out;
   MUX_Add12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg100_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg23_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg475_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg652_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg346_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg235_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg162_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg238_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg338_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg479_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg657_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg659_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg719_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg404_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg349_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg337_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg336_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_2_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_3_impl_out,
                 X => Delay1No58_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg248_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg248_out;
SharedReg310_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg312_out;
SharedReg491_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg557_out;
SharedReg657_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg657_out;
SharedReg555_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg555_out;
SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg683_out;
SharedReg736_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg736_out;
SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg362_out;
SharedReg730_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg730_out;
SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg425_out;
SharedReg554_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg554_out;
SharedReg644_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg644_out;
SharedReg311_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg311_out;
SharedReg113_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg113_out;
SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg362_out;
SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg11_out;
SharedReg7_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg7_out;
SharedReg365_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg365_out;
SharedReg552_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg552_out;
SharedReg486_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg486_out;
SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg425_out;
SharedReg109_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg109_out;
SharedReg169_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg169_out;
   MUX_Add12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg248_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg730_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg554_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg644_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg311_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg113_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg6_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg7_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg365_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg552_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg486_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg425_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg109_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg169_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg491_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg657_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg555_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg736_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg362_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_3_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_0_out,
                 Y => Delay1No58_out);

SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg348_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg348_out;
SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg362_out;
SharedReg490_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg490_out;
SharedReg642_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg642_out;
SharedReg668_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg668_out;
SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg637_out;
SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg552_out;
SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg729_out;
SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg482_out;
SharedReg738_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg738_out;
SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg729_out;
SharedReg420_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg420_out;
SharedReg313_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg313_out;
SharedReg363_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg363_out;
SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg362_out;
SharedReg111_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg111_out;
SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg482_out;
SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg27_out;
SharedReg23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg23_out;
SharedReg485_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg485_out;
SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg637_out;
SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg552_out;
SharedReg435_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg435_out;
SharedReg253_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg253_out;
SharedReg174_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg174_out;
   MUX_Add12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg738_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg420_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg313_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg363_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg111_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg22_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg362_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg485_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg435_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg253_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg174_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg490_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg642_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg668_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg637_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg552_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg729_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg482_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_3_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_4_impl_out,
                 X => Delay1No60_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg497_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg497_out;
SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg441_out;
SharedReg120_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg120_out;
SharedReg181_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg181_out;
SharedReg266_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg266_out;
SharedReg304_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg304_out;
SharedReg524_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg524_out;
SharedReg502_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg502_out;
SharedReg565_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg565_out;
SharedReg499_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg499_out;
SharedReg563_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg500_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg500_out;
SharedReg746_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg746_out;
SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg353_out;
SharedReg740_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg740_out;
SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg441_out;
SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg441_out;
SharedReg306_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg306_out;
SharedReg698_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg698_out;
SharedReg305_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg305_out;
SharedReg124_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg124_out;
SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg353_out;
SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg11_out;
SharedReg7_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg7_out;
SharedReg356_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg356_out;
   MUX_Add12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg497_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg499_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg500_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg746_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg740_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg306_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg698_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg441_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg305_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg124_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg353_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg6_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg7_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg356_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg120_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg181_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg266_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg304_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg524_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg502_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg565_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_4_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_0_out,
                 Y => Delay1No60_out);

SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg692_out;
SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg560_out;
SharedReg451_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg271_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg271_out;
SharedReg186_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg274_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg274_out;
SharedReg355_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg355_out;
SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg353_out;
SharedReg501_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg697_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg697_out;
SharedReg677_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg677_out;
SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg692_out;
SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg560_out;
SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg739_out;
SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg493_out;
SharedReg748_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg748_out;
SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg739_out;
SharedReg436_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg436_out;
SharedReg563_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg563_out;
SharedReg354_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg354_out;
SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg353_out;
SharedReg122_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg122_out;
SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg493_out;
SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg27_out;
SharedReg23_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg23_out;
SharedReg496_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg496_out;
   MUX_Add12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg677_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg692_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg560_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg748_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg739_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg436_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg563_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg354_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg451_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg122_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg493_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg22_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg23_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg496_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg271_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg186_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg274_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg355_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg353_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg697_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_4_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add121_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_0_impl_out,
                 X => Delay1No62_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast);

SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg538_out;
SharedReg15_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg8_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg539_out;
SharedReg752_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg752_out;
SharedReg542_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg542_out;
SharedReg192_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg192_out;
SharedReg704_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg704_out;
SharedReg773_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg773_out;
SharedReg507_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg507_out;
SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg539_out;
SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg749_out;
Delay17No20_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_15_cast <= Delay17No20_out;
SharedReg325_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg325_out;
SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg749_out;
SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg539_out;
SharedReg756_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg756_out;
SharedReg316_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg316_out;
SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg538_out;
SharedReg685_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg685_out;
SharedReg131_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg131_out;
SharedReg32_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg32_out;
SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg686_out;
SharedReg505_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg505_out;
SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg686_out;
SharedReg194_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg194_out;
   MUX_Add121_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg773_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg507_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay17No20_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg325_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg749_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg756_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg316_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg13_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg538_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg685_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg131_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg32_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg505_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg686_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg194_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg14_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg539_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg752_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg542_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg192_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg704_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_0_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_0_out,
                 Y => Delay1No62_out);

SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg685_out;
SharedReg31_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg30_out;
SharedReg24_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg686_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg686_out;
SharedReg689_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg689_out;
SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg749_out;
SharedReg200_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg200_out;
SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg579_out;
SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg579_out;
SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg541_out;
SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg685_out;
SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg541_out;
SharedReg544_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg544_out;
Delay43No_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_16_cast <= Delay43No_out;
SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg541_out;
SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg749_out;
SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg749_out;
SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg452_out;
SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg685_out;
SharedReg687_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg687_out;
SharedReg127_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg127_out;
SharedReg188_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg188_out;
SharedReg750_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg750_out;
SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg452_out;
SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg749_out;
SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg135_out;
   MUX_Add121_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg544_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay43No_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg541_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg29_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg685_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg687_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg127_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg188_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg750_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg452_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg30_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg686_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg689_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg749_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg200_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg579_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_0_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add121_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_1_impl_out,
                 X => Delay1No64_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast);

SharedReg143_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg40_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg646_out;
SharedReg514_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg514_out;
SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg646_out;
SharedReg212_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg212_out;
SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg545_out;
SharedReg15_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg14_out;
SharedReg8_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg546_out;
SharedReg662_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg662_out;
SharedReg549_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg549_out;
SharedReg210_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg210_out;
SharedReg714_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg714_out;
SharedReg785_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg785_out;
SharedReg516_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg516_out;
SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg546_out;
SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg659_out;
Delay17No21_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_21_cast <= Delay17No21_out;
SharedReg335_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg335_out;
SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg659_out;
SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg546_out;
SharedReg666_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg666_out;
SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg326_out;
SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg545_out;
SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg326_out;
   MUX_Add121_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg662_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg549_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg210_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg714_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg785_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg516_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay17No21_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg335_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg659_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg546_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg666_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg326_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg514_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg646_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg212_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg545_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg15_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg14_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_1_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_0_out,
                 Y => Delay1No64_out);

SharedReg139_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg139_out;
SharedReg206_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg206_out;
SharedReg660_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg660_out;
SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg462_out;
SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg659_out;
SharedReg147_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg645_out;
SharedReg31_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg30_out;
SharedReg24_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg646_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg646_out;
SharedReg649_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg649_out;
SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg659_out;
SharedReg218_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg218_out;
SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg593_out;
SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg593_out;
SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg548_out;
SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg645_out;
SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg548_out;
SharedReg551_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg551_out;
Delay43No1_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_22_cast <= Delay43No1_out;
SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg548_out;
SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg659_out;
SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg659_out;
SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg462_out;
SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg645_out;
SharedReg647_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg647_out;
   MUX_Add121_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg139_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg646_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg649_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg218_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg593_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg660_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg551_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay43No1_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg548_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg647_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg462_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg659_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg645_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg31_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg30_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_1_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add121_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_2_impl_out,
                 X => Delay1No66_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast);

SharedReg290_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg675_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg675_out;
SharedReg336_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg336_out;
SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg346_out;
SharedReg652_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg652_out;
SharedReg155_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg155_out;
SharedReg48_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg48_out;
SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg653_out;
SharedReg296_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg296_out;
SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg653_out;
SharedReg230_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg230_out;
SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg346_out;
SharedReg15_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg14_out;
SharedReg8_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg347_out;
SharedReg671_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg671_out;
SharedReg350_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg350_out;
SharedReg228_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg228_out;
SharedReg724_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg724_out;
SharedReg797_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg797_out;
SharedReg298_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg298_out;
SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg347_out;
SharedReg668_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg668_out;
Delay17No22_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_26_cast <= Delay17No22_out;
SharedReg345_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg345_out;
SharedReg472_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg472_out;
   MUX_Add121_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg675_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg230_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg15_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg13_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg14_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg671_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg350_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg228_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg336_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg724_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg797_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg298_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg347_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg668_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay17No22_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg345_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg472_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg346_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg652_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg155_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg48_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg296_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg653_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_2_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_2_impl_0_out,
                 Y => Delay1No66_out);

SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg668_out;
SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg668_out;
SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg472_out;
SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg652_out;
SharedReg654_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg654_out;
SharedReg151_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg151_out;
SharedReg224_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg224_out;
SharedReg669_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg669_out;
SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg472_out;
SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg668_out;
SharedReg159_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg652_out;
SharedReg31_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg30_out;
SharedReg24_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg24_out;
SharedReg653_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg653_out;
SharedReg656_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg656_out;
SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg668_out;
SharedReg236_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg236_out;
SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg607_out;
SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg607_out;
SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg349_out;
SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg652_out;
SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg349_out;
SharedReg352_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg352_out;
Delay43No2_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_27_cast <= Delay43No2_out;
SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg349_out;
   MUX_Add121_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg31_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg29_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg30_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg24_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg653_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg656_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg236_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg607_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg352_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay43No2_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg349_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg652_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg654_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg151_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg224_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg669_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg472_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg668_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_2_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_2_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add121_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_3_impl_out,
                 X => Delay1No68_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast);

SharedReg525_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg525_out;
SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg553_out;
SharedReg677_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg677_out;
Delay17No23_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast <= Delay17No23_out;
SharedReg371_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg371_out;
SharedReg482_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg482_out;
SharedReg311_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg311_out;
SharedReg489_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg489_out;
SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg362_out;
SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg552_out;
SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg362_out;
SharedReg167_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg167_out;
SharedReg56_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg56_out;
SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg638_out;
SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg523_out;
SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg638_out;
SharedReg248_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg248_out;
SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg552_out;
SharedReg15_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg14_out;
SharedReg8_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg8_out;
SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg553_out;
SharedReg680_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg680_out;
SharedReg556_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg556_out;
SharedReg246_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg246_out;
SharedReg734_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg734_out;
SharedReg809_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg809_out;
   MUX_Add121_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg525_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg167_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg56_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg638_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg248_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg15_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg13_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg677_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg14_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg8_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg553_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg680_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg556_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg246_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg734_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg809_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay17No23_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg371_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg482_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg311_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg489_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg362_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg552_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_3_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_0_out,
                 Y => Delay1No68_out);

SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg555_out;
SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg637_out;
SharedReg313_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg313_out;
SharedReg559_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg559_out;
Delay43No3_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast <= Delay43No3_out;
SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg555_out;
SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg677_out;
SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg677_out;
SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg482_out;
SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg637_out;
SharedReg639_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg639_out;
SharedReg163_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg163_out;
SharedReg242_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg242_out;
SharedReg678_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg678_out;
SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg482_out;
SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg677_out;
SharedReg171_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg171_out;
SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg637_out;
SharedReg31_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg30_out;
SharedReg24_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg24_out;
SharedReg638_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg638_out;
SharedReg641_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg641_out;
SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg677_out;
SharedReg254_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg254_out;
SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg621_out;
SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg621_out;
   MUX_Add121_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg639_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg163_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg242_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg678_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg171_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg31_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg29_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg313_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg30_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg24_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg638_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg641_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg254_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg621_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg559_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay43No3_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg555_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg677_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg482_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg637_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_3_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add121_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_4_impl_out,
                 X => Delay1No70_out_to_Add121_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add121_4_impl_parent_implementedSystem_port_1_cast);

SharedReg761_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg761_out;
SharedReg564_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg564_out;
SharedReg264_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg264_out;
SharedReg744_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg744_out;
SharedReg821_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg821_out;
SharedReg532_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg532_out;
SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg305_out;
SharedReg758_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg758_out;
Delay17No24_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast <= Delay17No24_out;
SharedReg361_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg361_out;
SharedReg493_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg493_out;
SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg305_out;
SharedReg765_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg765_out;
SharedReg353_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg353_out;
SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg560_out;
SharedReg692_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg692_out;
SharedReg179_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg179_out;
SharedReg64_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg64_out;
SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg693_out;
SharedReg531_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg531_out;
SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg693_out;
SharedReg266_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg266_out;
SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg14_out;
SharedReg8_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg8_out;
SharedReg561_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg561_out;
   MUX_Add121_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg761_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg564_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg493_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg765_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg353_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg692_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg179_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg64_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg531_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg264_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg693_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg266_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg560_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg15_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg13_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg14_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg8_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg561_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg744_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg821_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg532_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg305_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg758_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay17No24_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg361_out_to_MUX_Add121_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_4_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_4_impl_0_out,
                 Y => Delay1No70_out);

SharedReg696_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg696_out;
SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg758_out;
SharedReg272_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg272_out;
SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg635_out;
SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg635_out;
SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg692_out;
SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg563_out;
SharedReg566_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg566_out;
Delay43No4_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast <= Delay43No4_out;
SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg563_out;
SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg758_out;
SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg758_out;
SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg493_out;
SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg692_out;
SharedReg694_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg694_out;
SharedReg175_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg175_out;
SharedReg260_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg260_out;
SharedReg759_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg759_out;
SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg493_out;
SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg758_out;
SharedReg183_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg183_out;
SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg692_out;
SharedReg31_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg30_out;
SharedReg24_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg24_out;
SharedReg693_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg693_out;
   MUX_Add121_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg696_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg694_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg175_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg260_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg759_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg493_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg272_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg758_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg183_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg31_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg29_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg30_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg24_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg693_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg635_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg692_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg563_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg566_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay43No4_out_to_MUX_Add121_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add121_4_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_4_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No72_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg840_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg840_out;
SharedReg841_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg841_out;
SharedReg190_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg190_out;
SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg874_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg874_out;
SharedReg33_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg33_out;
SharedReg827_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg827_out;
SharedReg889_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg889_out;
SharedReg829_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg829_out;
SharedReg830_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg830_out;
SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg900_out;
SharedReg569_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg569_out;
SharedReg917_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg917_out;
SharedReg918_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg918_out;
SharedReg866_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg866_out;
SharedReg846_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg847_out;
SharedReg848_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg848_out;
SharedReg922_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg922_out;
SharedReg850_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg850_out;
SharedReg907_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg907_out;
SharedReg855_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg856_out;
SharedReg769_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg769_out;
SharedReg836_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg836_out;
SharedReg837_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg837_out;
SharedReg838_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg838_out;
SharedReg839_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg839_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg840_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg841_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg569_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg917_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg918_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg866_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg846_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg848_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg922_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg850_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg190_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg907_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg769_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg836_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg837_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg838_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg839_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg874_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg33_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg827_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg889_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg829_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg830_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No72_out);

SharedReg187_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg128_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg128_out;
SharedReg872_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg872_out;
SharedReg191_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg875_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg875_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg567_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg74_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg74_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg32_out;
SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg700_out;
SharedReg899_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg899_out;
SharedReg703_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg703_out;
SharedReg571_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg37_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg32_out;
SharedReg775_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg775_out;
SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg38_out;
SharedReg774_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg774_out;
SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg78_out;
SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg38_out;
SharedReg882_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg882_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg700_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg32_out;
SharedReg127_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg127_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg899_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg703_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg775_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg872_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg774_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg78_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg882_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg700_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg127_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg191_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg875_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg567_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg74_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No74_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg856_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg856_out;
SharedReg781_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg781_out;
SharedReg836_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg836_out;
SharedReg837_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg837_out;
SharedReg838_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg838_out;
SharedReg839_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg840_out;
SharedReg841_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg841_out;
SharedReg208_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg208_out;
SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg843_out;
SharedReg874_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg874_out;
SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg41_out;
SharedReg827_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg827_out;
SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg889_out;
SharedReg829_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg829_out;
SharedReg830_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg830_out;
SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg900_out;
SharedReg583_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg583_out;
SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg917_out;
SharedReg918_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg918_out;
SharedReg866_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg866_out;
SharedReg846_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg847_out;
SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg913_out;
SharedReg922_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg922_out;
SharedReg850_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg850_out;
SharedReg907_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg907_out;
SharedReg855_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg855_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg856_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg781_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg874_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg41_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg827_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg829_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg830_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg583_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg918_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg836_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg866_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg846_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg922_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg850_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg907_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg855_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg837_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg838_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg839_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg840_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg841_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg208_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No74_out);

SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg882_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg40_out;
SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg710_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg139_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg205_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg205_out;
SharedReg140_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg140_out;
SharedReg872_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg872_out;
SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg209_out;
SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg41_out;
SharedReg875_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg875_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg40_out;
SharedReg581_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg581_out;
SharedReg85_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg85_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg40_out;
SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg710_out;
SharedReg899_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg899_out;
SharedReg713_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg713_out;
SharedReg585_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg585_out;
SharedReg45_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg45_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg40_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg40_out;
SharedReg709_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg709_out;
SharedReg787_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg787_out;
SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg46_out;
SharedReg786_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg786_out;
SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg89_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg875_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg581_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg85_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg899_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg713_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg585_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg45_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg709_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg787_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg46_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg786_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg710_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg205_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg140_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg872_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No76_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg848_out;
SharedReg905_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg905_out;
SharedReg850_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg850_out;
SharedReg907_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg907_out;
SharedReg855_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg856_out;
SharedReg793_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg793_out;
SharedReg836_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg836_out;
SharedReg837_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg838_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg838_out;
SharedReg839_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg840_out;
SharedReg841_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg841_out;
SharedReg226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg226_out;
SharedReg843_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg843_out;
SharedReg874_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg874_out;
SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg49_out;
SharedReg827_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg827_out;
SharedReg889_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg889_out;
SharedReg829_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg829_out;
SharedReg830_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg830_out;
SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg900_out;
SharedReg597_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg597_out;
SharedReg833_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg833_out;
SharedReg918_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg918_out;
SharedReg866_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg866_out;
SharedReg846_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg847_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg905_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg839_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg840_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg841_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg843_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg874_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg827_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg889_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg829_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg850_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg830_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg597_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg833_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg918_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg866_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg846_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg847_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg907_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg856_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg793_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg836_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg838_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No76_out);

SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg792_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg798_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg798_out;
SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg882_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg882_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg720_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg48_out;
SharedReg151_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg223_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg223_out;
SharedReg152_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg152_out;
SharedReg872_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg872_out;
SharedReg227_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg227_out;
SharedReg49_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg49_out;
SharedReg875_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg875_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg48_out;
SharedReg595_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg595_out;
SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg96_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg48_out;
SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg720_out;
SharedReg899_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg899_out;
SharedReg154_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg154_out;
SharedReg599_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg599_out;
SharedReg53_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg53_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg48_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg223_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg152_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg872_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg227_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg49_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg875_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg595_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg899_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg154_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg599_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg53_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg798_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg882_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg720_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No78_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg917_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg917_out;
SharedReg880_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg880_out;
SharedReg854_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg49_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg49_out;
SharedReg848_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg848_out;
SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg94_out;
SharedReg852_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg852_out;
SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg94_out;
SharedReg891_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg891_out;
SharedReg871_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg871_out;
SharedReg842_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg842_out;
SharedReg843_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg843_out;
SharedReg901_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg901_out;
SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg853_out;
SharedReg791_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg791_out;
SharedReg828_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg828_out;
SharedReg153_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg153_out;
SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg225_out;
SharedReg406_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg406_out;
SharedReg899_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg899_out;
SharedReg827_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg827_out;
SharedReg154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg154_out;
SharedReg835_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg835_out;
SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg94_out;
SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg94_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg917_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg891_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg871_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg842_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg843_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg901_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg791_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg828_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg153_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg880_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg406_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg899_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg827_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg835_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg854_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg49_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg848_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg852_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No78_out);

SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg719_out;
SharedReg733_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg733_out;
SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg54_out;
SharedReg411_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg411_out;
SharedReg881_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg881_out;
SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg56_out;
SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg867_out;
SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg791_out;
SharedReg868_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg868_out;
SharedReg869_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg869_out;
SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg719_out;
SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg49_out;
SharedReg722_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg722_out;
SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg52_out;
SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg791_out;
SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg933_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg933_out;
SharedReg48_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg48_out;
SharedReg860_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg860_out;
SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg861_out;
SharedReg908_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg908_out;
SharedReg723_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg723_out;
SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg56_out;
SharedReg865_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg865_out;
SharedReg97_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg97_out;
SharedReg876_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg877_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg733_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg869_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg719_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg722_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg933_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg48_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg860_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg908_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg723_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg865_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg97_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg876_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg411_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg881_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg56_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg791_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg868_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No80_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg827_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg827_out;
SharedReg828_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg829_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg829_out;
SharedReg830_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg830_out;
SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg625_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg625_out;
SharedReg833_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg833_out;
SharedReg918_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg918_out;
SharedReg866_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg866_out;
SharedReg846_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg847_out;
SharedReg848_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg848_out;
SharedReg905_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg905_out;
SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg850_out;
SharedReg907_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg907_out;
SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg856_out;
SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg817_out;
SharedReg836_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg836_out;
SharedReg837_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg837_out;
SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg838_out;
SharedReg839_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg840_out;
SharedReg117_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg117_out;
SharedReg262_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg262_out;
SharedReg843_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg843_out;
SharedReg874_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg874_out;
SharedReg65_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg65_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg827_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg848_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg905_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg907_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg856_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg836_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg837_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg829_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg839_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg840_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg117_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg262_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg843_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg874_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg65_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg830_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg625_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg833_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg918_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg866_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg846_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No80_out);

SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg64_out;
SharedReg116_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg116_out;
SharedReg118_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg740_out;
SharedReg899_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg899_out;
SharedReg178_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg627_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg627_out;
SharedReg69_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg69_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg64_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg64_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg64_out;
SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg70_out;
SharedReg822_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg822_out;
SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg122_out;
SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg70_out;
SharedReg882_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg882_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg64_out;
SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg740_out;
SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg64_out;
SharedReg175_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg175_out;
SharedReg259_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg259_out;
SharedReg871_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg871_out;
SharedReg872_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg872_out;
SharedReg263_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg263_out;
SharedReg65_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg875_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg875_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg822_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg882_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg118_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg175_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg259_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg871_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg872_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg263_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg875_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg740_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg627_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg69_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg64_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product11_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_3_impl_out,
                 X => Delay1No82_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg611_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg611_out;
SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg833_out;
SharedReg918_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg866_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg866_out;
SharedReg846_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg847_out;
SharedReg913_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg913_out;
SharedReg922_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg922_out;
SharedReg850_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg907_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg907_out;
SharedReg855_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg856_out;
SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg805_out;
SharedReg836_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg836_out;
SharedReg837_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg837_out;
SharedReg838_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg838_out;
SharedReg839_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg840_out;
SharedReg841_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg841_out;
SharedReg244_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg244_out;
SharedReg843_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg843_out;
SharedReg874_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg874_out;
SharedReg57_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg57_out;
SharedReg858_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg858_out;
SharedReg889_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg889_out;
SharedReg829_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg829_out;
SharedReg830_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg830_out;
SharedReg900_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg900_out;
   MUX_Product11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg611_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg856_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg836_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg837_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg838_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg839_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg840_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg841_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg244_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg843_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg874_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg57_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg858_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg889_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg829_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg830_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg900_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg866_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg846_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg913_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg922_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg907_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_3_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_0_out,
                 Y => Delay1No82_out);

SharedReg899_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg166_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg166_out;
SharedReg613_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg613_out;
SharedReg61_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg61_out;
SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg56_out;
SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg56_out;
SharedReg729_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg729_out;
SharedReg811_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg811_out;
SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg62_out;
SharedReg810_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg810_out;
SharedReg111_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg111_out;
SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg62_out;
SharedReg882_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg882_out;
SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg56_out;
SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg730_out;
SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg56_out;
SharedReg163_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg163_out;
SharedReg241_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg241_out;
SharedReg164_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg164_out;
SharedReg872_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg872_out;
SharedReg245_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg245_out;
SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg57_out;
SharedReg875_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg875_out;
SharedReg420_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg420_out;
SharedReg609_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg609_out;
SharedReg107_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg107_out;
SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg56_out;
SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg730_out;
   MUX_Product11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg111_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg882_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg163_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg241_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg164_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg872_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg613_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg245_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg875_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg420_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg609_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg730_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg61_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg56_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg729_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg811_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg62_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg810_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_3_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No84_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg870_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg870_out;
SharedReg841_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg841_out;
SharedReg893_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg893_out;
SharedReg843_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg844_out;
SharedReg845_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg845_out;
SharedReg858_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg921_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg921_out;
SharedReg74_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg74_out;
SharedReg894_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg894_out;
SharedReg900_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg900_out;
SharedReg898_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg898_out;
SharedReg703_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg703_out;
SharedReg920_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg920_out;
SharedReg927_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg927_out;
SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg847_out;
SharedReg878_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg878_out;
SharedReg849_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg916_out;
SharedReg855_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg887_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg887_out;
SharedReg857_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg857_out;
SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg836_out;
SharedReg852_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg838_out;
SharedReg869_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg869_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg870_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg841_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg900_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg898_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg703_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg920_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg927_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg847_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg878_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg849_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg880_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg893_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg916_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg887_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg857_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg852_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg838_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg869_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg845_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg921_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg74_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg894_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No84_out);

SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg569_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg33_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg33_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg767_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg767_out;
SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg860_out;
SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg703_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg703_out;
SharedReg919_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg919_out;
SharedReg571_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg772_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg72_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg72_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg32_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg72_out;
SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg38_out;
SharedReg774_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg774_out;
SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg38_out;
SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg38_out;
SharedReg577_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg577_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg72_out;
SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg128_out;
SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg72_out;
SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg127_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg703_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg919_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg774_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg38_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg577_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg72_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg127_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg767_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No86_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg887_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg887_out;
SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg857_out;
SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg836_out;
SharedReg852_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg838_out;
SharedReg869_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg869_out;
SharedReg870_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg870_out;
SharedReg841_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg841_out;
SharedReg893_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg893_out;
SharedReg843_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg843_out;
SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg844_out;
SharedReg845_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg845_out;
SharedReg858_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg858_out;
SharedReg921_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg921_out;
SharedReg85_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg85_out;
SharedReg894_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg894_out;
SharedReg900_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg900_out;
SharedReg898_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg898_out;
SharedReg713_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg713_out;
SharedReg920_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg920_out;
SharedReg927_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg927_out;
SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg847_out;
SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg904_out;
SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg916_out;
SharedReg855_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg855_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg887_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg845_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg858_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg921_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg85_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg894_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg900_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg898_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg713_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg920_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg927_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg847_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg880_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg916_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg855_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg838_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg870_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg841_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg893_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg843_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No86_out);

SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg591_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg591_out;
SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg140_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg139_out;
SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg583_out;
SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg41_out;
SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg41_out;
SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg41_out;
SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg40_out;
SharedReg779_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg779_out;
SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg860_out;
SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg390_out;
SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg390_out;
SharedReg713_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg713_out;
SharedReg919_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg919_out;
SharedReg585_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg585_out;
SharedReg784_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg784_out;
SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg83_out;
SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg83_out;
SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg583_out;
SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg83_out;
SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg46_out;
SharedReg786_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg786_out;
SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg46_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg591_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg779_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg390_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg713_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg919_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg585_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg784_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg786_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg46_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg140_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg139_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg583_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No88_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg878_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg878_out;
SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg880_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg855_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg887_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg887_out;
SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg857_out;
SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg836_out;
SharedReg852_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg838_out;
SharedReg869_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg869_out;
SharedReg870_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg870_out;
SharedReg841_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg841_out;
SharedReg893_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg893_out;
SharedReg843_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg843_out;
SharedReg844_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg844_out;
SharedReg845_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg845_out;
SharedReg858_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg858_out;
SharedReg921_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg921_out;
SharedReg96_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg96_out;
SharedReg894_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg894_out;
SharedReg900_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg900_out;
SharedReg898_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg898_out;
SharedReg154_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg154_out;
SharedReg920_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg920_out;
SharedReg927_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg927_out;
SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg847_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg878_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg869_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg870_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg841_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg893_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg843_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg844_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg845_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg858_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg921_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg96_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg880_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg894_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg900_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg898_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg154_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg920_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg927_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg847_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg887_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg852_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg838_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No88_out);

SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg914_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg914_out;
SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg798_out;
SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg54_out;
SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg605_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg605_out;
SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg94_out;
SharedReg152_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg152_out;
SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg151_out;
SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg49_out;
SharedReg597_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg597_out;
SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg49_out;
SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg49_out;
SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg49_out;
SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg48_out;
SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg791_out;
SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg860_out;
SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg406_out;
SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg406_out;
SharedReg723_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg723_out;
SharedReg864_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg864_out;
SharedReg599_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg599_out;
SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg796_out;
SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg94_out;
SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg94_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg914_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg151_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg597_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg49_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg406_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg723_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg864_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg599_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg605_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg152_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No90_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg733_out;
SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg54_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg54_out;
SharedReg886_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg851_out;
SharedReg878_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg878_out;
SharedReg836_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg836_out;
SharedReg883_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg883_out;
SharedReg923_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg923_out;
SharedReg924_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg924_out;
SharedReg891_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg891_out;
SharedReg95_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg95_out;
SharedReg842_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg842_out;
SharedReg873_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg873_out;
SharedReg909_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg909_out;
SharedReg853_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg853_out;
SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg858_out;
SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg828_out;
SharedReg890_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg890_out;
SharedReg861_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg861_out;
SharedReg831_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg832_out;
SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg858_out;
SharedReg834_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg834_out;
SharedReg866_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg866_out;
SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg903_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg924_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg891_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg95_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg842_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg873_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg909_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg853_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg890_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg861_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg831_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg832_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg858_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg834_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg866_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg54_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg886_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg878_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg836_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg883_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg923_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No90_out);

SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg719_out;
SharedReg919_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg919_out;
SharedReg720_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg720_out;
SharedReg885_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg411_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg411_out;
SharedReg792_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg792_out;
SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg56_out;
SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg791_out;
SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg791_out;
SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg719_out;
SharedReg595_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg595_out;
SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg791_out;
SharedReg871_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg871_out;
SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg794_out;
SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg52_out;
SharedReg721_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg721_out;
SharedReg152_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg152_out;
SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg404_out;
SharedReg94_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg94_out;
SharedReg405_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg405_out;
SharedReg224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg224_out;
SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg50_out;
SharedReg154_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg154_out;
SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg56_out;
SharedReg227_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg227_out;
SharedReg97_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg97_out;
SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg404_out;
SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg719_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg919_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg595_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg871_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg721_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg152_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg94_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg405_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg720_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg154_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg227_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg97_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg404_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg885_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg411_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg792_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg56_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg719_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product21_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_4_impl_out,
                 X => Delay1No92_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast);

SharedReg858_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg858_out;
SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg116_out;
SharedReg118_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg894_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg894_out;
SharedReg900_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg898_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg898_out;
SharedReg178_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg920_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg920_out;
SharedReg927_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg927_out;
SharedReg846_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg847_out;
SharedReg878_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg878_out;
SharedReg816_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg880_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg916_out;
SharedReg855_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg855_out;
SharedReg887_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg887_out;
SharedReg857_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg857_out;
SharedReg836_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg836_out;
SharedReg852_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg838_out;
SharedReg869_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg869_out;
SharedReg870_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg870_out;
SharedReg892_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg892_out;
SharedReg893_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg893_out;
SharedReg843_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg843_out;
SharedReg844_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg844_out;
SharedReg845_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg845_out;
   MUX_Product21_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg858_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg847_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg878_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg880_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg916_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg855_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg887_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg857_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg836_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg852_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg118_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg838_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg869_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg870_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg892_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg893_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg843_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg844_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg845_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg894_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg898_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg920_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg927_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg846_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_4_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_0_out,
                 Y => Delay1No92_out);

SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg64_out;
SharedReg859_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg859_out;
SharedReg860_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg860_out;
SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg438_out;
SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg438_out;
SharedReg743_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg743_out;
SharedReg864_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg864_out;
SharedReg627_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg627_out;
SharedReg820_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg820_out;
SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg116_out;
SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg64_out;
SharedReg914_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg914_out;
SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg70_out;
SharedReg822_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg822_out;
SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg70_out;
SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg70_out;
SharedReg633_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg633_out;
SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg116_out;
SharedReg176_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg176_out;
SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg116_out;
SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg175_out;
SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg175_out;
SharedReg437_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg437_out;
SharedReg625_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg625_out;
SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg65_out;
SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg65_out;
   MUX_Product21_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg859_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg64_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg914_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg822_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg70_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg633_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg176_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg860_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg437_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg625_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg65_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg438_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg743_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg864_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg627_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg820_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_4_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product31_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_3_impl_out,
                 X => Delay1No94_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast);

SharedReg898_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg898_out;
SharedReg166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg166_out;
SharedReg920_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg927_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg927_out;
SharedReg846_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg846_out;
SharedReg847_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg847_out;
SharedReg904_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg904_out;
SharedReg849_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg916_out;
SharedReg855_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg887_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg887_out;
SharedReg857_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg857_out;
SharedReg836_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg836_out;
SharedReg852_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg838_out;
SharedReg869_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg869_out;
SharedReg870_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg870_out;
SharedReg841_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg841_out;
SharedReg893_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg893_out;
SharedReg843_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg843_out;
SharedReg844_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg844_out;
SharedReg845_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg845_out;
SharedReg609_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg609_out;
SharedReg921_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg921_out;
SharedReg107_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg107_out;
SharedReg894_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg894_out;
SharedReg900_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg900_out;
   MUX_Product31_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg898_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg887_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg857_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg836_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg852_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg838_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg869_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg870_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg841_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg893_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg843_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg844_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg845_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg609_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg921_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg894_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg900_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg927_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg846_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg847_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg904_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg849_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg880_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg916_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product31_3_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_0_out,
                 Y => Delay1No94_out);

SharedReg733_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg864_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg864_out;
SharedReg613_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg613_out;
SharedReg808_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg105_out;
SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg611_out;
SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg62_out;
SharedReg810_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg810_out;
SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg62_out;
SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg62_out;
SharedReg619_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg619_out;
SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg105_out;
SharedReg164_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg164_out;
SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg105_out;
SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg163_out;
SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg163_out;
SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg57_out;
SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg611_out;
SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg57_out;
SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg57_out;
SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg57_out;
SharedReg858_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg858_out;
SharedReg803_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg803_out;
SharedReg860_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg860_out;
SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg422_out;
   MUX_Product31_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg864_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg619_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg164_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg163_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg613_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg57_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg858_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg803_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg860_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg422_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg808_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg611_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg62_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg810_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product31_3_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No96_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg277_out;
SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg280_out;
SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg282_out;
SharedReg386_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg386_out;
SharedReg384_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg384_out;
SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg567_out;
SharedReg504_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg504_out;
SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg279_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg277_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg277_out;
SharedReg316_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg316_out;
SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg452_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg277_out;
SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg452_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg277_out;
SharedReg128_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg277_out;
SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg567_out;
SharedReg699_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg699_out;
SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg279_out;
SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg279_out;
SharedReg317_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg317_out;
SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg573_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg504_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg316_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg452_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg699_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg279_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg317_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg386_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg384_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No96_out);

SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg453_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg453_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg277_out;
SharedReg755_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg755_out;
SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg378_out;
SharedReg573_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg573_out;
SharedReg699_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg699_out;
SharedReg685_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg685_out;
SharedReg316_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg316_out;
SharedReg505_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg505_out;
SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg504_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg277_out;
SharedReg510_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg510_out;
SharedReg317_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg317_out;
SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg687_out;
SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg504_out;
SharedReg82_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg82_out;
SharedReg452_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg452_out;
SharedReg769_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg769_out;
SharedReg373_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg373_out;
SharedReg459_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg459_out;
SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg461_out;
SharedReg540_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg540_out;
SharedReg385_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg385_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg699_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg685_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg316_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg505_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg510_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg317_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg504_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg82_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg452_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg769_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg373_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg459_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg540_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg385_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg453_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg277_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg755_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg573_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No98_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg709_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg709_out;
SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg285_out;
SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg285_out;
SharedReg327_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg327_out;
SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg587_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg283_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg283_out;
SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg286_out;
SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg288_out;
SharedReg402_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg402_out;
SharedReg400_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg400_out;
SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg581_out;
SharedReg513_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg513_out;
SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg285_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg283_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg283_out;
SharedReg326_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg326_out;
SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg462_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg283_out;
SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg462_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg283_out;
SharedReg140_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg140_out;
SharedReg504_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg504_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg709_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg402_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg400_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg581_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg513_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg326_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg462_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg140_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg504_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg285_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg327_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg283_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No98_out);

SharedReg781_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg781_out;
SharedReg389_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg469_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg471_out;
SharedReg547_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg401_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg401_out;
SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg513_out;
SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg463_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg283_out;
SharedReg665_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg665_out;
SharedReg394_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg394_out;
SharedReg587_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg587_out;
SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg709_out;
SharedReg645_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg645_out;
SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg326_out;
SharedReg514_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg514_out;
SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg513_out;
SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg283_out;
SharedReg519_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg519_out;
SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg327_out;
SharedReg647_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg647_out;
SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg513_out;
SharedReg93_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg93_out;
SharedReg685_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg685_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg781_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg665_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg394_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg587_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg645_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg514_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg469_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg283_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg519_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg647_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg93_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg685_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg401_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No100_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg289_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg472_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg289_out;
SharedReg152_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg289_out;
SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg719_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg719_out;
SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg515_out;
SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg291_out;
SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg337_out;
SharedReg601_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg601_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg289_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg2_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg289_out;
SharedReg292_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg292_out;
SharedReg294_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg294_out;
SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg418_out;
SharedReg416_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg416_out;
SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg595_out;
SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg295_out;
SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg291_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg289_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg289_out;
SharedReg336_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg336_out;
SharedReg645_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg645_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg601_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg292_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg294_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg416_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg336_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg645_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg152_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg719_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg291_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No100_out);

SharedReg546_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg546_out;
SharedReg338_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg295_out;
SharedReg104_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg104_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg472_out;
SharedReg793_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg793_out;
SharedReg405_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
SharedReg479_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg479_out;
SharedReg481_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg481_out;
SharedReg348_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg348_out;
SharedReg417_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg417_out;
SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg295_out;
SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg18_out;
SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg473_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg289_out;
SharedReg674_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg674_out;
SharedReg410_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg410_out;
SharedReg601_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg601_out;
SharedReg719_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg719_out;
SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg652_out;
SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg336_out;
SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg296_out;
SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg295_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg289_out;
SharedReg301_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg301_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg546_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg417_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg674_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg410_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg601_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg719_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg295_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg301_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg104_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg793_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg479_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg481_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg348_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No102_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg522_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg522_out;
SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg297_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg310_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg310_out;
SharedReg362_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg362_out;
SharedReg652_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg652_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg310_out;
SharedReg482_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg482_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg310_out;
SharedReg164_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg164_out;
SharedReg295_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg295_out;
SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg609_out;
SharedReg729_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg729_out;
SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg312_out;
SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg312_out;
SharedReg363_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg363_out;
SharedReg615_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg615_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg310_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg2_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg310_out;
SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg313_out;
SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg315_out;
SharedReg434_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg434_out;
SharedReg432_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg432_out;
SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg609_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg522_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg295_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg729_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg363_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg615_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg434_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg432_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg609_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg362_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg652_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg482_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg164_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No102_out);

SharedReg637_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg637_out;
SharedReg362_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg362_out;
SharedReg523_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg523_out;
SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg522_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg310_out;
SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg673_out;
SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg347_out;
SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg364_out;
SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg522_out;
SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg115_out;
SharedReg652_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg652_out;
SharedReg805_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg805_out;
SharedReg421_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg421_out;
SharedReg490_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg490_out;
SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg492_out;
SharedReg554_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg554_out;
SharedReg433_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg433_out;
SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg522_out;
SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg18_out;
SharedReg483_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg483_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg310_out;
SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg683_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg426_out;
SharedReg615_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg615_out;
SharedReg729_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg729_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg637_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg362_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg652_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg805_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg421_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg490_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg554_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg433_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg523_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg483_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg615_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg729_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg522_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No104_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg307_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg307_out;
SharedReg309_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg309_out;
SharedReg450_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg450_out;
SharedReg448_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg448_out;
SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg623_out;
SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg677_out;
SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg306_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg304_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg304_out;
SharedReg353_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg353_out;
SharedReg637_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg637_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg304_out;
SharedReg493_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg493_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg304_out;
SharedReg176_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg176_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg304_out;
SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg623_out;
SharedReg739_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg739_out;
SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg524_out;
SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg306_out;
SharedReg354_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg354_out;
SharedReg629_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg629_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg304_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg9_out;
SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg2_out;
SharedReg522_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg522_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg309_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg637_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg493_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg176_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg739_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg450_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg354_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg629_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg522_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg448_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg623_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg306_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg353_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No104_out);

SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg764_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg764_out;
SharedReg442_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg442_out;
SharedReg629_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg629_out;
SharedReg739_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg739_out;
SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg353_out;
SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg353_out;
SharedReg531_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg531_out;
SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg530_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg304_out;
SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg535_out;
SharedReg553_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg553_out;
SharedReg355_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg355_out;
SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg530_out;
SharedReg126_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg126_out;
SharedReg493_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg493_out;
SharedReg817_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg817_out;
SharedReg437_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg437_out;
SharedReg643_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg643_out;
SharedReg503_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg503_out;
SharedReg562_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg562_out;
SharedReg449_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg449_out;
SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg530_out;
SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg18_out;
SharedReg494_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg494_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg764_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg553_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg355_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg126_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg493_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg817_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg437_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg643_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg503_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg442_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg562_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg449_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg494_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg629_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg353_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg531_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg304_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product12_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_0_impl_out,
                 X => Delay1No106_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg187_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg841_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg841_out;
SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg33_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg33_out;
SharedReg901_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg901_out;
SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg768_out;
SharedReg931_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg931_out;
SharedReg767_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg767_out;
SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg829_out;
SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg569_out;
SharedReg908_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg908_out;
SharedReg898_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg898_out;
SharedReg932_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg932_out;
SharedReg834_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg834_out;
SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg835_out;
SharedReg876_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg877_out;
SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg72_out;
SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg72_out;
SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg850_out;
SharedReg77_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg77_out;
SharedReg886_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg851_out;
SharedReg577_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg577_out;
SharedReg867_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg867_out;
SharedReg883_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg883_out;
SharedReg868_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg868_out;
SharedReg839_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg839_out;
   MUX_Product12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg841_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg908_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg898_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg932_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg834_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg876_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg877_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg72_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg77_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg886_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg851_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg577_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg867_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg883_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg868_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg839_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg33_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg901_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg931_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg767_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg569_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_0_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_0_out,
                 Y => Delay1No106_out);

SharedReg870_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg870_out;
SharedReg73_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg897_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg897_out;
SharedReg873_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg873_out;
SharedReg701_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg701_out;
SharedReg910_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg910_out;
SharedReg767_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg767_out;
SharedReg926_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg926_out;
SharedReg129_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg129_out;
SharedReg894_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg894_out;
SharedReg700_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg700_out;
SharedReg569_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg569_out;
SharedReg771_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg771_out;
SharedReg130_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg130_out;
SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg76_out;
SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg32_out;
SharedReg878_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg878_out;
SharedReg879_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg879_out;
SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg33_out;
SharedReg885_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg885_out;
SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg38_out;
SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg33_out;
SharedReg888_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg888_out;
SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg128_out;
SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg32_out;
SharedReg72_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg72_out;
   MUX_Product12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg870_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg700_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg569_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg771_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg130_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg878_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg879_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg897_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg885_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg33_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg888_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg72_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg873_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg701_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg910_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg767_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg926_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg129_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg894_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_0_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product12_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_1_impl_out,
                 X => Delay1No108_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg851_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg851_out;
SharedReg591_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg591_out;
SharedReg867_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg867_out;
SharedReg883_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg868_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg868_out;
SharedReg839_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg839_out;
SharedReg205_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg205_out;
SharedReg841_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg841_out;
SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg583_out;
SharedReg41_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg41_out;
SharedReg901_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg901_out;
SharedReg780_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg780_out;
SharedReg931_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg931_out;
SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg779_out;
SharedReg829_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg829_out;
SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg583_out;
SharedReg908_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg908_out;
SharedReg898_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg898_out;
SharedReg932_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg932_out;
SharedReg834_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg834_out;
SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg835_out;
SharedReg876_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg877_out;
SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg904_out;
SharedReg83_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg83_out;
SharedReg850_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg850_out;
SharedReg88_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg88_out;
SharedReg886_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg886_out;
   MUX_Product12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg851_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg591_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg901_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg780_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg931_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg829_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg908_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg898_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg932_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg834_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg867_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg876_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg877_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg83_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg850_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg88_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg886_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg883_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg868_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg839_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg205_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg841_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg583_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg41_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_1_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_0_out,
                 Y => Delay1No108_out);

SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg888_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg888_out;
SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg40_out;
SharedReg140_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg83_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg83_out;
SharedReg870_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg870_out;
SharedReg84_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg84_out;
SharedReg897_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg897_out;
SharedReg873_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg873_out;
SharedReg711_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg711_out;
SharedReg910_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg910_out;
SharedReg779_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg926_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg926_out;
SharedReg141_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg141_out;
SharedReg894_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg894_out;
SharedReg710_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg710_out;
SharedReg583_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg583_out;
SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg783_out;
SharedReg142_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg142_out;
SharedReg87_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg87_out;
SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg40_out;
SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg40_out;
SharedReg582_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg582_out;
SharedReg879_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg879_out;
SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg41_out;
SharedReg885_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg885_out;
SharedReg46_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg46_out;
   MUX_Product12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg888_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg711_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg910_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg926_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg141_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg894_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg710_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg583_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg142_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg87_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg582_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg879_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg41_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg885_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg46_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg140_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg83_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg870_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg84_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg897_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg873_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_1_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product12_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_2_impl_out,
                 X => Delay1No110_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg94_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg596_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg850_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg850_out;
SharedReg99_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg886_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg851_out;
SharedReg605_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg605_out;
SharedReg867_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg867_out;
SharedReg883_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg883_out;
SharedReg868_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg868_out;
SharedReg839_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg839_out;
SharedReg223_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg223_out;
SharedReg841_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg841_out;
SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg597_out;
SharedReg49_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg49_out;
SharedReg901_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg901_out;
SharedReg792_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg792_out;
SharedReg931_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg931_out;
SharedReg791_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg791_out;
SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg829_out;
SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg597_out;
SharedReg908_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg908_out;
SharedReg898_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg898_out;
SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg834_out;
SharedReg835_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg835_out;
SharedReg876_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg877_out;
   MUX_Product12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg839_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg223_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg841_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg49_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg901_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg792_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg931_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg791_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg850_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg597_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg908_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg898_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg834_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg835_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg876_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg877_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg99_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg886_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg851_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg605_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg867_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg883_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg868_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_2_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_0_out,
                 Y => Delay1No110_out);

SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg878_out;
SharedReg914_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg914_out;
SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg49_out;
SharedReg885_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg54_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg54_out;
SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg49_out;
SharedReg888_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg888_out;
SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg152_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg152_out;
SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg48_out;
SharedReg94_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg94_out;
SharedReg870_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg870_out;
SharedReg95_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg95_out;
SharedReg897_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg897_out;
SharedReg873_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg873_out;
SharedReg721_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg721_out;
SharedReg910_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg910_out;
SharedReg791_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg791_out;
SharedReg926_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg926_out;
SharedReg153_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg153_out;
SharedReg894_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg894_out;
SharedReg720_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg720_out;
SharedReg597_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg597_out;
SharedReg228_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg228_out;
SharedReg154_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg154_out;
SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg98_out;
SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg48_out;
   MUX_Product12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg914_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg94_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg870_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg95_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg897_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg873_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg721_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg910_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg791_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg926_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg153_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg894_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg720_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg597_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg228_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg154_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg885_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg54_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg49_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg888_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg152_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_2_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product12_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_3_impl_out,
                 X => Delay1No112_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg898_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg898_out;
SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg834_out;
SharedReg835_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg835_out;
SharedReg876_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg877_out;
SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg904_out;
SharedReg105_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg850_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg110_out;
SharedReg886_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg851_out;
SharedReg619_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg619_out;
SharedReg867_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg867_out;
SharedReg883_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg883_out;
SharedReg868_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg868_out;
SharedReg839_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg839_out;
SharedReg241_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg241_out;
SharedReg841_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg841_out;
SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg611_out;
SharedReg57_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg57_out;
SharedReg901_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg901_out;
SharedReg804_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg804_out;
SharedReg935_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg935_out;
SharedReg803_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg803_out;
SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg829_out;
SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg611_out;
SharedReg908_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg908_out;
   MUX_Product12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg898_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg886_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg851_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg619_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg867_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg883_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg868_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg839_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg241_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg841_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg834_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg57_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg901_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg804_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg935_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg803_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg611_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg908_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg835_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg876_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg877_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_3_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_0_out,
                 Y => Delay1No112_out);

SharedReg611_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg611_out;
SharedReg246_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg246_out;
SharedReg166_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg166_out;
SharedReg109_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg109_out;
SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg56_out;
SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg56_out;
SharedReg610_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg610_out;
SharedReg879_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg879_out;
SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg57_out;
SharedReg885_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg885_out;
SharedReg62_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg62_out;
SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg57_out;
SharedReg888_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg888_out;
SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg56_out;
SharedReg164_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg164_out;
SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg56_out;
SharedReg105_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg105_out;
SharedReg870_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg870_out;
SharedReg106_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg106_out;
SharedReg897_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg897_out;
SharedReg873_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg873_out;
SharedReg731_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg731_out;
SharedReg910_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg910_out;
SharedReg729_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg729_out;
SharedReg926_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg926_out;
SharedReg165_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg165_out;
SharedReg894_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg894_out;
SharedReg730_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg730_out;
   MUX_Product12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg611_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg246_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg62_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg888_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg164_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg105_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg870_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg106_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg897_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg166_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg873_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg731_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg910_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg729_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg926_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg165_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg894_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg730_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg109_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg56_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg610_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg879_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg57_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg885_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_3_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product12_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_4_impl_out,
                 X => Delay1No114_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg931_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg931_out;
SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg829_out;
SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg625_out;
SharedReg908_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg898_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg898_out;
SharedReg833_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg834_out;
SharedReg835_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg835_out;
SharedReg876_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg877_out;
SharedReg116_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg116_out;
SharedReg624_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg624_out;
SharedReg850_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg850_out;
SharedReg121_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg121_out;
SharedReg886_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg851_out;
SharedReg633_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg633_out;
SharedReg867_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg867_out;
SharedReg883_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg883_out;
SharedReg868_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg868_out;
SharedReg839_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg839_out;
SharedReg259_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg259_out;
SharedReg896_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg896_out;
SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg625_out;
SharedReg65_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg65_out;
SharedReg901_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg901_out;
SharedReg816_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg816_out;
   MUX_Product12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg931_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg877_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg116_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg624_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg850_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg121_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg886_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg633_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg867_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg883_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg868_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg839_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg259_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg896_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg65_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg901_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg816_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg625_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg898_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg833_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg834_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg835_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg876_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_4_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_0_out,
                 Y => Delay1No114_out);

SharedReg815_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg815_out;
SharedReg259_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg259_out;
SharedReg177_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg177_out;
SharedReg894_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg894_out;
SharedReg740_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg740_out;
SharedReg625_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg625_out;
SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg264_out;
SharedReg178_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg178_out;
SharedReg120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg120_out;
SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg64_out;
SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg64_out;
SharedReg878_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg878_out;
SharedReg914_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg914_out;
SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg65_out;
SharedReg885_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg885_out;
SharedReg70_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg70_out;
SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg65_out;
SharedReg888_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg888_out;
SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg64_out;
SharedReg176_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg176_out;
SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg64_out;
SharedReg116_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg116_out;
SharedReg870_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg870_out;
SharedReg437_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg437_out;
SharedReg897_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg897_out;
SharedReg873_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg873_out;
SharedReg741_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg741_out;
SharedReg910_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg910_out;
   MUX_Product12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg815_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg259_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg878_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg914_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg885_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg70_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg65_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg888_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg176_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg177_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg116_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg870_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg437_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg897_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg873_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg741_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg910_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg894_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg740_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg625_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg178_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg64_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_4_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No116_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg891_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg891_out;
SharedReg871_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg871_out;
SharedReg842_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg842_out;
SharedReg843_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg901_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg901_out;
SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg853_out;
SharedReg767_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg767_out;
SharedReg828_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg828_out;
SharedReg129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg129_out;
SharedReg189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg189_out;
SharedReg374_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg899_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg899_out;
SharedReg934_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg934_out;
SharedReg130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg130_out;
SharedReg835_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg835_out;
SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg72_out;
SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg72_out;
SharedReg904_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg904_out;
SharedReg849_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg880_out;
SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg33_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg33_out;
SharedReg848_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg848_out;
SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg72_out;
SharedReg852_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg852_out;
SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg72_out;
SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg72_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg891_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg871_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg899_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg934_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg835_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg904_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg849_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg880_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg842_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg33_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg848_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg852_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg72_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg901_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg767_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg828_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No116_out);

SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg702_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg767_out;
SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg73_out;
SharedReg933_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg933_out;
SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg32_out;
SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg860_out;
SharedReg861_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg861_out;
SharedReg908_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg908_out;
SharedReg703_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg703_out;
SharedReg771_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg771_out;
SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg865_out;
SharedReg75_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg75_out;
SharedReg876_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg877_out;
SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg699_out;
SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg73_out;
SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg33_out;
SharedReg38_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg38_out;
SharedReg379_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg379_out;
SharedReg881_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg881_out;
SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg40_out;
SharedReg867_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg867_out;
SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg767_out;
SharedReg868_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg868_out;
SharedReg869_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg869_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg908_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg703_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg771_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg75_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg876_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg877_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg699_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg702_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg38_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg379_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg881_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg867_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg868_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg869_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg767_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg73_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg933_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg861_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No118_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg41_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg922_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg922_out;
SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg852_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg83_out;
SharedReg891_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg891_out;
SharedReg871_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg871_out;
SharedReg842_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg842_out;
SharedReg843_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg843_out;
SharedReg901_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg901_out;
SharedReg853_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg853_out;
SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg828_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg828_out;
SharedReg141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg141_out;
SharedReg207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg207_out;
SharedReg390_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg390_out;
SharedReg899_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg899_out;
SharedReg934_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg934_out;
SharedReg142_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg142_out;
SharedReg835_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg835_out;
SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg83_out;
SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg83_out;
SharedReg917_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg917_out;
SharedReg849_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg880_out;
SharedReg854_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg855_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg922_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg901_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg853_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg828_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg390_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg899_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg934_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg142_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg835_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg917_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg849_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg880_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg854_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg855_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg83_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg891_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg871_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg842_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg843_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No118_out);

SharedReg881_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg881_out;
SharedReg799_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg867_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg867_out;
SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg779_out;
SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg868_out;
SharedReg869_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg869_out;
SharedReg709_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg709_out;
SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg712_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg712_out;
SharedReg44_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg44_out;
SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg779_out;
SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg84_out;
SharedReg933_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg933_out;
SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg40_out;
SharedReg860_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg860_out;
SharedReg861_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg861_out;
SharedReg908_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg908_out;
SharedReg713_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg713_out;
SharedReg783_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg783_out;
SharedReg865_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg865_out;
SharedReg86_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg86_out;
SharedReg876_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg877_out;
SharedReg723_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg723_out;
SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg84_out;
SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg41_out;
SharedReg46_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg46_out;
SharedReg395_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg395_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg881_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg933_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg860_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg861_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg908_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg713_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg783_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg865_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg867_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg86_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg876_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg877_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg723_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg84_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg46_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg395_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg779_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg709_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg712_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg44_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No120_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg889_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg889_out;
SharedReg166_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg166_out;
SharedReg835_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg835_out;
SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg105_out;
SharedReg917_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg917_out;
SharedReg849_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg849_out;
SharedReg880_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg880_out;
SharedReg854_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg57_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg57_out;
SharedReg922_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg922_out;
SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg105_out;
SharedReg852_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg852_out;
SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg105_out;
SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg105_out;
SharedReg891_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg891_out;
SharedReg871_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg871_out;
SharedReg842_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg842_out;
SharedReg843_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg843_out;
SharedReg901_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg901_out;
SharedReg853_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg853_out;
SharedReg841_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg841_out;
SharedReg828_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg828_out;
SharedReg165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg165_out;
SharedReg243_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg243_out;
SharedReg422_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg422_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg889_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg57_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg922_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg852_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg891_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg871_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg842_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg166_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg843_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg901_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg853_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg841_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg828_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg243_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg422_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg835_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg105_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg917_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg849_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg880_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg854_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No120_out);

SharedReg733_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg623_out;
SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg865_out;
SharedReg108_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg108_out;
SharedReg876_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg877_out;
SharedReg743_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg743_out;
SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg106_out;
SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg57_out;
SharedReg62_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg427_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg427_out;
SharedReg881_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg881_out;
SharedReg823_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg823_out;
SharedReg867_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg867_out;
SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg803_out;
SharedReg868_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg868_out;
SharedReg869_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg869_out;
SharedReg729_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg729_out;
SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg57_out;
SharedReg732_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg732_out;
SharedReg60_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg60_out;
SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg803_out;
SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg106_out;
SharedReg176_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg176_out;
SharedReg56_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg56_out;
SharedReg860_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg860_out;
SharedReg861_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg861_out;
SharedReg908_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg908_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg427_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg881_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg823_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg867_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg868_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg869_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg729_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg732_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg60_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg803_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg176_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg56_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg860_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg861_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg908_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg108_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg876_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg877_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg743_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg106_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No122_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg177_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg116_out;
SharedReg65_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg65_out;
SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg116_out;
SharedReg178_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg178_out;
SharedReg261_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
SharedReg438_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg438_out;
SharedReg815_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg815_out;
SharedReg899_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg899_out;
SharedReg843_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg843_out;
SharedReg842_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg842_out;
SharedReg891_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg891_out;
SharedReg901_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg901_out;
SharedReg853_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg853_out;
SharedReg880_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg880_out;
SharedReg904_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg904_out;
SharedReg852_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg852_out;
SharedReg854_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg835_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg835_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg815_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg899_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg843_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg842_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg891_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg901_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg853_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg880_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg904_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg852_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg854_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg835_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg65_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg178_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg438_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product32_4_impl_0_LUT_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No122_out);

SharedReg68_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg117_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg70_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg119_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg119_out;
SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg815_out;
SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg815_out;
SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg739_out;
SharedReg443_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg443_out;
SharedReg743_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg743_out;
SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg860_out;
SharedReg742_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg742_out;
SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg739_out;
SharedReg908_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg908_out;
SharedReg933_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg933_out;
SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg867_out;
SharedReg868_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg868_out;
SharedReg869_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg869_out;
SharedReg865_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg865_out;
SharedReg881_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg881_out;
SharedReg876_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg876_out;
SharedReg877_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg877_out;
SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg861_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg742_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg908_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg933_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg868_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg869_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg865_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg881_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg876_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg877_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg70_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg119_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg815_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg739_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg443_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg743_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product32_4_impl_1_LUT_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No124_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg891_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg891_out;
SharedReg73_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg842_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg842_out;
SharedReg873_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg873_out;
SharedReg909_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg909_out;
SharedReg853_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg853_out;
SharedReg858_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg828_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg828_out;
SharedReg890_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg890_out;
SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg861_out;
SharedReg831_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg832_out;
SharedReg833_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg834_out;
SharedReg866_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg866_out;
SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg903_out;
SharedReg913_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg913_out;
SharedReg905_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg905_out;
SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg906_out;
SharedReg38_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg38_out;
SharedReg886_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg851_out;
SharedReg878_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg878_out;
SharedReg836_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg836_out;
SharedReg883_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg883_out;
SharedReg923_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg923_out;
SharedReg924_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg924_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg891_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg831_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg832_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg833_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg834_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg866_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg913_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg905_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg842_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg38_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg886_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg851_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg878_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg836_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg883_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg923_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg924_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg873_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg909_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg853_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg828_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg890_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No124_out);

SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg871_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg871_out;
SharedReg770_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg770_out;
SharedReg36_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg701_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg701_out;
SharedReg128_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg128_out;
SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg372_out;
SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg72_out;
SharedReg373_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg373_out;
SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg34_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg34_out;
SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg130_out;
SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg130_out;
SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg191_out;
SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg75_out;
SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg372_out;
SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg699_out;
SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg699_out;
SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg768_out;
SharedReg700_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg700_out;
SharedReg885_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg885_out;
SharedReg379_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg379_out;
SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg768_out;
SharedReg40_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg40_out;
SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg767_out;
SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg767_out;
SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg699_out;
SharedReg567_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg567_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg871_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg34_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg130_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg700_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg770_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg885_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg379_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg768_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg40_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg699_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg567_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg701_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg372_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg373_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product6_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_1_impl_out,
                 X => Delay1No126_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg851_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg851_out;
SharedReg849_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg849_out;
SharedReg836_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg836_out;
SharedReg883_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg923_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg923_out;
SharedReg924_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg924_out;
SharedReg891_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg891_out;
SharedReg84_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg84_out;
SharedReg842_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg842_out;
SharedReg873_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg873_out;
SharedReg909_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg909_out;
SharedReg853_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg853_out;
SharedReg858_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg858_out;
SharedReg828_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg828_out;
SharedReg890_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg890_out;
SharedReg861_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg861_out;
SharedReg831_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg832_out;
SharedReg833_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg834_out;
SharedReg866_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg866_out;
SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg903_out;
SharedReg723_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg723_out;
SharedReg905_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg905_out;
SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg906_out;
SharedReg46_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg46_out;
SharedReg886_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg886_out;
   MUX_Product6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg851_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg849_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg909_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg853_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg858_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg828_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg890_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg861_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg831_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg832_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg833_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg834_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg836_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg866_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg723_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg905_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg46_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg886_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg883_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg923_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg924_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg891_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg84_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg842_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg873_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_1_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_0_out,
                 Y => Delay1No126_out);

SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg780_out;
SharedReg94_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg779_out;
SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg779_out;
SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg709_out;
SharedReg581_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg581_out;
SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg779_out;
SharedReg871_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg871_out;
SharedReg782_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg782_out;
SharedReg44_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg44_out;
SharedReg711_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg711_out;
SharedReg140_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg140_out;
SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg388_out;
SharedReg83_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg83_out;
SharedReg389_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg389_out;
SharedReg206_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg206_out;
SharedReg42_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg42_out;
SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg142_out;
SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg142_out;
SharedReg209_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg209_out;
SharedReg86_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg86_out;
SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg388_out;
SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg709_out;
SharedReg919_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg919_out;
SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg780_out;
SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg710_out;
SharedReg885_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg885_out;
SharedReg395_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg395_out;
   MUX_Product6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg711_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg140_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg83_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg389_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg206_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg42_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg142_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg209_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg86_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg388_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg919_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg780_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg885_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg395_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg709_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg581_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg779_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg871_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg782_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg44_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_1_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product6_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_3_impl_out,
                 X => Delay1No128_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast);

SharedReg832_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg832_out;
SharedReg921_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg921_out;
SharedReg834_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg834_out;
SharedReg866_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg866_out;
SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
SharedReg743_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg743_out;
SharedReg905_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg905_out;
SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg906_out;
SharedReg62_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg886_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg886_out;
SharedReg851_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg851_out;
SharedReg849_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg849_out;
SharedReg836_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg836_out;
SharedReg883_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg883_out;
SharedReg923_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg923_out;
SharedReg924_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg924_out;
SharedReg891_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg891_out;
SharedReg106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg106_out;
SharedReg842_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg842_out;
SharedReg873_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg873_out;
SharedReg909_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg909_out;
SharedReg853_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg853_out;
SharedReg841_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg841_out;
SharedReg828_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg828_out;
SharedReg890_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg890_out;
SharedReg861_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg861_out;
SharedReg831_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg831_out;
   MUX_Product6_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg832_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg921_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg886_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg851_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg849_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg836_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg883_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg923_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg924_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg891_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg842_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg834_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg873_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg909_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg853_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg841_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg828_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg890_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg861_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg831_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg866_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg743_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg905_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_3_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_0_out,
                 Y => Delay1No128_out);

SharedReg166_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg815_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg815_out;
SharedReg245_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg108_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg108_out;
SharedReg420_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg420_out;
SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg729_out;
SharedReg919_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg919_out;
SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg804_out;
SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg730_out;
SharedReg885_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg885_out;
SharedReg427_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg427_out;
SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg804_out;
SharedReg116_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg116_out;
SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg803_out;
SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg803_out;
SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg729_out;
SharedReg609_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg609_out;
SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg803_out;
SharedReg871_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg871_out;
SharedReg806_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg806_out;
SharedReg60_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg60_out;
SharedReg731_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg731_out;
SharedReg164_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg164_out;
SharedReg65_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg65_out;
SharedReg105_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg105_out;
SharedReg421_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg421_out;
SharedReg242_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg242_out;
SharedReg58_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg58_out;
   MUX_Product6_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg815_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg427_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg116_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg609_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg803_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg871_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg806_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg245_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg60_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg731_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg164_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg65_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg105_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg421_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg242_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg58_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg108_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg420_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg729_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg919_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg804_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg885_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_3_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product6_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_4_impl_out,
                 X => Delay1No130_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg70_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg890_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg890_out;
SharedReg924_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg924_out;
SharedReg836_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg836_out;
SharedReg873_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg873_out;
SharedReg842_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg842_out;
SharedReg891_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg891_out;
SharedReg923_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg923_out;
SharedReg832_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg832_out;
SharedReg909_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg909_out;
SharedReg853_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg853_out;
SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg906_out;
SharedReg913_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg913_out;
SharedReg851_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg851_out;
SharedReg883_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg883_out;
SharedReg834_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg834_out;
SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg831_out;
SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg902_out;
SharedReg886_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg886_out;
SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg903_out;
SharedReg866_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg866_out;
SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg861_out;
SharedReg858_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg858_out;
   MUX_Product6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg890_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg853_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg913_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg851_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg883_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg834_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg886_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg924_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg866_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg858_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg836_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg873_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg842_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg891_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg923_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg832_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg909_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product6_4_impl_0_LUT_out,
                 oMux => MUX_Product6_4_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_0_out,
                 Y => Delay1No130_out);

SharedReg68_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg178_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg178_out;
SharedReg263_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg263_out;
SharedReg66_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg66_out;
SharedReg119_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg119_out;
SharedReg260_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg260_out;
SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg436_out;
SharedReg741_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg741_out;
SharedReg623_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg623_out;
SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg815_out;
SharedReg437_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg437_out;
SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg739_out;
SharedReg740_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg740_out;
SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg815_out;
SharedReg816_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg816_out;
SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg739_out;
SharedReg443_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg443_out;
SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg436_out;
SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg739_out;
SharedReg818_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg818_out;
SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg815_out;
SharedReg885_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg885_out;
   MUX_Product6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg437_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg740_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg816_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg443_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg739_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg178_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg818_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg815_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg885_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg263_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg66_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg119_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg260_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg436_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg741_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg623_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product6_4_impl_1_LUT_out,
                 oMux => MUX_Product6_4_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Subtract4_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_0_impl_out,
                 X => Delay1No132_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg316_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg316_out;
SharedReg686_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg686_out;
SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg504_out;
SharedReg137_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg137_out;
SharedReg193_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg193_out;
SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg72_out;
SharedReg567_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg34_out;
SharedReg539_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg539_out;
SharedReg322_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg322_out;
SharedReg324_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg324_out;
SharedReg511_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg511_out;
SharedReg540_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg540_out;
SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg504_out;
SharedReg538_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg538_out;
SharedReg277_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg277_out;
SharedReg749_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg749_out;
SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg72_out;
SharedReg187_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg187_out;
SharedReg453_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg453_out;
SharedReg278_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg278_out;
SharedReg505_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg505_out;
SharedReg705_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg705_out;
   MUX_Subtract4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg539_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg322_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg324_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg511_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg540_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg538_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg277_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg749_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg72_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg187_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg453_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg278_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg505_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg705_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg10_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg316_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg686_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg504_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg137_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg193_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_0_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_0_out,
                 Y => Delay1No132_out);

SharedReg79_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg538_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg538_out;
SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg452_out;
SharedReg508_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg508_out;
SharedReg76_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg76_out;
SharedReg201_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg201_out;
SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg767_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg767_out;
SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg127_out;
SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg452_out;
SharedReg281_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg281_out;
Delay18No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast <= Delay18No15_out;
SharedReg755_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg755_out;
SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg504_out;
SharedReg509_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg509_out;
SharedReg749_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg749_out;
SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg504_out;
SharedReg750_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg750_out;
SharedReg188_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg188_out;
SharedReg33_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg33_out;
SharedReg454_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg454_out;
SharedReg757_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg757_out;
SharedReg751_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg751_out;
Delay27No10_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast <= Delay27No10_out;
   MUX_Subtract4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg767_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg127_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg281_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay18No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg755_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg509_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg749_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg750_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg188_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg33_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg454_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg757_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg751_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay27No10_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg26_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg538_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg452_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg508_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg76_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg201_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_0_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No134_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg205_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg463_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg463_out;
SharedReg284_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg284_out;
SharedReg514_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg514_out;
SharedReg715_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg715_out;
SharedReg92_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg92_out;
SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg326_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg326_out;
SharedReg646_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg646_out;
SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg513_out;
SharedReg149_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg149_out;
SharedReg211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg211_out;
SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg83_out;
SharedReg581_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg581_out;
SharedReg42_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg42_out;
SharedReg546_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg546_out;
SharedReg332_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg332_out;
SharedReg334_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg334_out;
SharedReg520_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg520_out;
SharedReg547_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg547_out;
SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg513_out;
SharedReg545_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg545_out;
SharedReg283_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg283_out;
SharedReg462_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg462_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg326_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg646_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg149_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg83_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg581_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg42_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg546_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg463_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg332_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg334_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg520_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg547_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg513_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg545_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg283_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg462_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg284_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg514_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg715_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg92_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg10_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No134_out);

SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg41_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg464_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg464_out;
SharedReg667_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg667_out;
SharedReg661_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg661_out;
Delay27No11_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= Delay27No11_out;
SharedReg90_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg90_out;
SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg26_out;
SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg545_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg545_out;
SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg462_out;
SharedReg517_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg517_out;
SharedReg87_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg87_out;
SharedReg219_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg219_out;
SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg139_out;
SharedReg779_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg779_out;
SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg139_out;
SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg462_out;
SharedReg287_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg287_out;
Delay18No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast <= Delay18No16_out;
SharedReg665_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg665_out;
SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg513_out;
SharedReg518_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg518_out;
SharedReg659_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg659_out;
SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg513_out;
SharedReg660_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg660_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg545_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg517_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg87_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg219_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg779_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg139_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg462_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg464_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg287_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay18No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg665_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg518_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg659_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg513_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg660_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg667_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay27No11_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg90_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg26_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Subtract4_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_2_impl_out,
                 X => Delay1No136_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg348_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg295_out;
SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg289_out;
SharedReg668_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg668_out;
SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg223_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg223_out;
SharedReg473_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg473_out;
SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg290_out;
SharedReg296_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg296_out;
SharedReg725_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg725_out;
SharedReg103_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg103_out;
SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg7_out;
SharedReg336_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg336_out;
SharedReg653_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg653_out;
SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg295_out;
SharedReg161_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg161_out;
SharedReg229_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg229_out;
SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg94_out;
SharedReg595_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg595_out;
SharedReg50_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg50_out;
SharedReg347_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg347_out;
SharedReg342_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg342_out;
SharedReg344_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg344_out;
SharedReg302_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg302_out;
   MUX_Subtract4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg725_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg103_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg10_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg336_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg653_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg295_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg161_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg229_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg595_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg50_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg347_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg342_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg344_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg302_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg668_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg223_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg473_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg296_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_2_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_0_out,
                 Y => Delay1No136_out);

SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg295_out;
SharedReg300_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg668_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg668_out;
SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg295_out;
SharedReg669_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg669_out;
SharedReg224_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg224_out;
SharedReg49_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg49_out;
SharedReg647_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg647_out;
SharedReg676_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg676_out;
SharedReg670_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg670_out;
Delay27No12_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast <= Delay27No12_out;
SharedReg101_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg101_out;
SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg26_out;
SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg23_out;
SharedReg346_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg346_out;
SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg472_out;
SharedReg299_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg299_out;
SharedReg98_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg98_out;
SharedReg237_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg237_out;
SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg151_out;
SharedReg791_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg791_out;
SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg151_out;
SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg472_out;
SharedReg293_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg293_out;
Delay18No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast <= Delay18No17_out;
SharedReg674_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg674_out;
   MUX_Subtract4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay27No12_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg101_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg26_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg346_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg299_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg98_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg668_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg237_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg791_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg151_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg472_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg293_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay18No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg674_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg295_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg669_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg224_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg49_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg647_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg676_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg670_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_2_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Subtract4_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_3_impl_out,
                 X => Delay1No138_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg609_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg58_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg58_out;
SharedReg553_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg368_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg368_out;
SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg370_out;
SharedReg528_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg528_out;
SharedReg554_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg522_out;
SharedReg552_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg552_out;
SharedReg310_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg310_out;
SharedReg482_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg482_out;
SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg105_out;
SharedReg241_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg241_out;
SharedReg483_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg483_out;
SharedReg311_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg311_out;
SharedReg523_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg523_out;
SharedReg735_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg735_out;
SharedReg114_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg114_out;
SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg7_out;
SharedReg362_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg362_out;
SharedReg638_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg638_out;
SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg522_out;
SharedReg173_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg173_out;
SharedReg247_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg247_out;
SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg105_out;
   MUX_Subtract4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg482_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg241_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg483_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg311_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg523_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg735_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg114_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg553_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg10_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg362_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg638_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg173_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg247_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg105_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg368_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg528_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg522_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg552_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg310_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_3_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_0_out,
                 Y => Delay1No138_out);

SharedReg803_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg163_out;
SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg482_out;
SharedReg314_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg314_out;
Delay18No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast <= Delay18No18_out;
SharedReg683_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg683_out;
SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg522_out;
SharedReg527_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg527_out;
SharedReg677_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg677_out;
SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg522_out;
SharedReg678_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg678_out;
SharedReg242_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg242_out;
SharedReg57_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg57_out;
SharedReg484_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg484_out;
SharedReg684_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg684_out;
SharedReg679_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg679_out;
Delay27No13_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast <= Delay27No13_out;
SharedReg112_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg112_out;
SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg26_out;
SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg23_out;
SharedReg552_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg552_out;
SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg482_out;
SharedReg526_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg526_out;
SharedReg109_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg109_out;
SharedReg255_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg255_out;
SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg163_out;
   MUX_Subtract4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg678_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg242_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg57_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg484_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg684_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg679_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay27No13_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg112_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg26_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg552_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg526_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg109_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg255_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg163_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg314_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay18No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg683_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg527_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg677_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg522_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_3_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Subtract4_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_4_impl_out,
                 X => Delay1No140_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg354_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg354_out;
SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg530_out;
SharedReg185_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg185_out;
SharedReg265_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
SharedReg623_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg623_out;
SharedReg66_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg66_out;
SharedReg561_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg561_out;
SharedReg359_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg359_out;
SharedReg360_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg360_out;
SharedReg536_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg536_out;
SharedReg562_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg562_out;
SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg530_out;
SharedReg560_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg560_out;
SharedReg304_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg304_out;
SharedReg758_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg758_out;
SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg116_out;
SharedReg259_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg259_out;
SharedReg494_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg494_out;
SharedReg305_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg305_out;
SharedReg531_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg531_out;
SharedReg745_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg745_out;
SharedReg125_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg125_out;
SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg7_out;
SharedReg552_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg552_out;
   MUX_Subtract4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg354_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg536_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg562_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg530_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg560_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg304_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg758_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg259_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg494_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg305_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg185_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg531_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg745_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg125_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg10_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg552_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg265_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg623_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg66_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg561_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg359_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg360_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_4_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_0_out,
                 Y => Delay1No140_out);

SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg493_out;
SharedReg533_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg533_out;
SharedReg120_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg273_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg273_out;
SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg815_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg815_out;
SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg175_out;
SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg493_out;
SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg308_out;
Delay18No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast <= Delay18No19_out;
SharedReg764_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg764_out;
SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg530_out;
SharedReg534_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg534_out;
SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg758_out;
SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg530_out;
SharedReg759_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg759_out;
SharedReg260_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg260_out;
SharedReg65_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg65_out;
SharedReg639_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg639_out;
SharedReg766_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg766_out;
SharedReg760_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg760_out;
Delay27No14_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast <= Delay27No14_out;
SharedReg123_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg123_out;
SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg26_out;
SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg23_out;
SharedReg304_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg304_out;
   MUX_Subtract4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg533_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg764_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg534_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg530_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg759_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg260_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg65_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg639_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg766_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg120_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg760_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay27No14_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg123_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg26_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg304_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg273_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg815_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg175_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg493_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay18No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_4_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product37_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_4_impl_out,
                 X => Delay1No142_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast);

SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg863_out;
SharedReg815_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg815_out;
SharedReg865_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg865_out;
SharedReg936_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg936_out;
SharedReg911_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg912_out;
SharedReg932_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg932_out;
SharedReg804_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg804_out;
SharedReg906_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg906_out;
SharedReg854_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg856_out;
SharedReg116_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg116_out;
SharedReg867_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg867_out;
SharedReg852_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg852_out;
SharedReg928_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg928_out;
SharedReg609_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg609_out;
SharedReg895_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg895_out;
SharedReg892_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg892_out;
SharedReg872_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg872_out;
SharedReg925_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg925_out;
SharedReg901_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg901_out;
SharedReg884_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg884_out;
SharedReg841_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg841_out;
SharedReg105_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg105_out;
SharedReg860_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg860_out;
SharedReg244_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg244_out;
SharedReg58_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg58_out;
   MUX_Product37_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg815_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg116_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg867_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg852_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg928_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg609_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg895_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg892_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg872_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg865_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg925_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg901_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg884_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg841_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg105_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg860_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg244_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg58_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg936_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg911_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg932_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg804_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg906_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg854_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product37_4_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_0_out,
                 Y => Delay1No142_out);

SharedReg166_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg926_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg926_out;
SharedReg245_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg425_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg425_out;
SharedReg420_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg420_out;
SharedReg609_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg609_out;
SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg819_out;
SharedReg914_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg914_out;
SharedReg611_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg611_out;
SharedReg615_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg615_out;
SharedReg736_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg736_out;
SharedReg427_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg427_out;
SharedReg879_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg879_out;
SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg729_out;
SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg729_out;
SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg729_out;
SharedReg929_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg929_out;
SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg729_out;
SharedReg421_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg421_out;
SharedReg732_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg732_out;
SharedReg424_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg424_out;
SharedReg805_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg805_out;
SharedReg106_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg106_out;
SharedReg117_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg117_out;
SharedReg859_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg859_out;
SharedReg57_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg57_out;
SharedReg861_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg861_out;
SharedReg862_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg862_out;
   MUX_Product37_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg736_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg427_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg879_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg929_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg729_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg421_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg732_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg245_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg424_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg805_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg106_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg117_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg859_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg57_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg861_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg862_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg425_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg420_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg609_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg914_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg611_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg615_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product37_4_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Product18_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_2_impl_out,
                 X => Delay1No144_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg856_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg856_out;
SharedReg94_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg94_out;
SharedReg867_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg867_out;
SharedReg852_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg928_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg928_out;
SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg581_out;
SharedReg895_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg895_out;
SharedReg892_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg892_out;
SharedReg872_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg872_out;
SharedReg925_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg925_out;
SharedReg901_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg901_out;
SharedReg884_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg884_out;
SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg581_out;
SharedReg83_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg83_out;
SharedReg860_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg860_out;
SharedReg208_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg208_out;
SharedReg42_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg42_out;
SharedReg863_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg863_out;
SharedReg142_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg142_out;
SharedReg865_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg865_out;
SharedReg936_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg936_out;
SharedReg911_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg912_out;
SharedReg932_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg932_out;
SharedReg780_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg780_out;
SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg906_out;
SharedReg854_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg855_out;
   MUX_Product18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg856_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg901_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg884_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg83_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg860_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg208_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg42_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg863_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg142_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg865_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg867_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg936_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg911_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg912_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg932_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg780_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg854_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg855_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg928_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg581_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg895_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg892_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg872_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg925_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product18_2_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_0_out,
                 Y => Delay1No144_out);

SharedReg395_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg395_out;
SharedReg879_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg879_out;
SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg709_out;
SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg709_out;
SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg709_out;
SharedReg929_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg929_out;
SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg709_out;
SharedReg389_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg389_out;
SharedReg712_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg712_out;
SharedReg392_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg392_out;
SharedReg781_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg781_out;
SharedReg84_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg84_out;
SharedReg858_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg858_out;
SharedReg859_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg859_out;
SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg41_out;
SharedReg861_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg861_out;
SharedReg862_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg862_out;
SharedReg142_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg142_out;
SharedReg864_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg864_out;
SharedReg209_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg209_out;
SharedReg393_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg393_out;
SharedReg388_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg388_out;
SharedReg581_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg581_out;
SharedReg795_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg795_out;
SharedReg914_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg914_out;
SharedReg583_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg583_out;
SharedReg587_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg587_out;
SharedReg716_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg716_out;
   MUX_Product18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg395_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg879_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg781_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg858_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg859_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg861_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg862_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg142_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg864_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg209_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg393_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg388_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg581_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg795_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg914_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg583_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg587_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg716_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg709_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg389_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg712_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg392_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product18_2_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product18_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_3_impl_out,
                 X => Delay1No146_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg932_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg932_out;
SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg854_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg856_out;
SharedReg105_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg105_out;
SharedReg867_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg867_out;
SharedReg852_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg852_out;
SharedReg928_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg928_out;
SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg595_out;
SharedReg895_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg895_out;
SharedReg892_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg892_out;
SharedReg872_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg872_out;
SharedReg925_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg925_out;
SharedReg901_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg901_out;
SharedReg884_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg884_out;
SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg595_out;
SharedReg94_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg94_out;
SharedReg860_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg860_out;
SharedReg226_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg226_out;
SharedReg50_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg50_out;
SharedReg863_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg863_out;
SharedReg931_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg931_out;
SharedReg865_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg865_out;
SharedReg936_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg936_out;
SharedReg911_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg912_out;
   MUX_Product18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg932_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg895_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg892_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg872_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg925_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg901_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg884_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg595_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg94_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg860_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg226_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg50_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg863_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg931_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg865_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg936_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg911_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg912_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg854_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg856_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg105_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg867_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg852_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg928_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product18_3_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_0_out,
                 Y => Delay1No146_out);

SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg597_out;
SharedReg807_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg597_out;
SharedReg601_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg601_out;
SharedReg726_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg726_out;
SharedReg411_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg411_out;
SharedReg878_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg878_out;
SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg719_out;
SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg719_out;
SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg719_out;
SharedReg929_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg929_out;
SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg719_out;
SharedReg405_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg405_out;
SharedReg722_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg722_out;
SharedReg408_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg408_out;
SharedReg793_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg793_out;
SharedReg95_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg858_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg858_out;
SharedReg859_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg859_out;
SharedReg49_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg49_out;
SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg861_out;
SharedReg862_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg862_out;
SharedReg154_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg154_out;
SharedReg803_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg803_out;
SharedReg227_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg227_out;
SharedReg409_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg409_out;
SharedReg404_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg404_out;
SharedReg595_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg595_out;
   MUX_Product18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg929_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg405_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg722_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg408_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg793_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg858_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg859_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg49_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg597_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg862_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg154_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg803_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg227_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg409_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg404_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg595_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg601_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg726_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg411_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg878_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg719_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product18_3_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product28_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_2_impl_out,
                 X => Delay1No148_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast);

SharedReg887_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg887_out;
SharedReg849_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg849_out;
SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg779_out;
SharedReg883_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg924_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg924_out;
SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg779_out;
SharedReg896_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg896_out;
SharedReg782_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg782_out;
SharedReg930_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg930_out;
SharedReg781_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg781_out;
SharedReg140_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg140_out;
SharedReg935_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg935_out;
SharedReg828_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg828_out;
SharedReg711_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg711_out;
SharedReg830_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg830_out;
SharedReg831_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg832_out;
SharedReg833_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg833_out;
SharedReg865_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg865_out;
SharedReg938_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg938_out;
SharedReg581_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg581_out;
SharedReg709_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg709_out;
SharedReg934_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg934_out;
SharedReg582_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg582_out;
SharedReg915_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg915_out;
SharedReg587_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg587_out;
SharedReg716_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg716_out;
   MUX_Product28_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg887_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg849_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg781_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg140_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg935_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg828_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg711_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg830_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg831_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg832_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg833_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg865_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg938_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg581_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg709_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg934_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg582_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg915_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg587_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg716_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg883_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg924_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg779_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg896_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg782_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg930_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_2_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_0_out,
                 Y => Delay1No148_out);

SharedReg395_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg395_out;
SharedReg95_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg867_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg867_out;
SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg709_out;
SharedReg928_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg928_out;
SharedReg780_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg780_out;
SharedReg895_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg895_out;
SharedReg389_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg389_out;
SharedReg872_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg872_out;
SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg392_out;
SharedReg909_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg909_out;
SharedReg884_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg884_out;
SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg709_out;
SharedReg205_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg205_out;
SharedReg937_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg937_out;
SharedReg584_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg584_out;
SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg392_out;
SharedReg208_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg208_out;
SharedReg210_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg210_out;
SharedReg86_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg86_out;
SharedReg393_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg393_out;
SharedReg911_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg912_out;
SharedReg795_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg795_out;
SharedReg914_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg914_out;
SharedReg710_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg710_out;
SharedReg885_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg886_out;
   MUX_Product28_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg395_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg909_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg884_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg205_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg937_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg584_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg208_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg210_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg86_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg867_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg393_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg911_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg912_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg795_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg914_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg710_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg885_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg886_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg709_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg928_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg780_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg895_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg389_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg872_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg392_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_2_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product28_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_3_impl_out,
                 X => Delay1No150_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg934_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg915_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg915_out;
SharedReg601_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg601_out;
SharedReg726_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg726_out;
SharedReg887_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg887_out;
SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg904_out;
SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg791_out;
SharedReg883_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg883_out;
SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg791_out;
SharedReg924_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg924_out;
SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg791_out;
SharedReg896_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg896_out;
SharedReg794_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg794_out;
SharedReg930_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg930_out;
SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg793_out;
SharedReg152_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg152_out;
SharedReg935_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg935_out;
SharedReg828_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg828_out;
SharedReg721_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg721_out;
SharedReg830_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg830_out;
SharedReg831_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg832_out;
SharedReg803_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg803_out;
SharedReg865_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg865_out;
SharedReg938_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg938_out;
SharedReg595_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg595_out;
SharedReg719_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg719_out;
   MUX_Product28_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg924_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg896_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg794_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg930_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg152_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg935_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg828_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg721_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg915_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg830_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg831_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg832_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg803_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg865_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg938_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg595_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg719_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg601_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg726_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg887_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg904_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg883_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg791_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_3_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_0_out,
                 Y => Delay1No150_out);

SharedReg596_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg596_out;
SharedReg807_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg720_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg720_out;
SharedReg885_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg886_out;
SharedReg411_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg411_out;
SharedReg729_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg729_out;
SharedReg867_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg867_out;
SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg719_out;
SharedReg928_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg928_out;
SharedReg792_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg792_out;
SharedReg895_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg895_out;
SharedReg405_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg405_out;
SharedReg872_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg872_out;
SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg408_out;
SharedReg909_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg909_out;
SharedReg884_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg884_out;
SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg719_out;
SharedReg223_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg223_out;
SharedReg937_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg937_out;
SharedReg598_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg598_out;
SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg408_out;
SharedReg226_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg226_out;
SharedReg933_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg933_out;
SharedReg97_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg97_out;
SharedReg409_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg409_out;
SharedReg911_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg912_out;
   MUX_Product28_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg596_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg792_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg895_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg405_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg872_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg909_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg884_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg223_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg937_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg720_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg598_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg408_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg226_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg933_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg97_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg409_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg911_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg912_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg885_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg886_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg411_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg729_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg867_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg719_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg928_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_3_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product28_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_4_impl_out,
                 X => Delay1No152_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast);

SharedReg832_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg832_out;
SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg865_out;
SharedReg938_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg938_out;
SharedReg609_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg609_out;
SharedReg729_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg729_out;
SharedReg934_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg934_out;
SharedReg610_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg610_out;
SharedReg915_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg915_out;
SharedReg615_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg615_out;
SharedReg736_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg736_out;
SharedReg887_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg887_out;
SharedReg849_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg849_out;
SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg803_out;
SharedReg883_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg883_out;
SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg803_out;
SharedReg924_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg924_out;
SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg803_out;
SharedReg896_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg896_out;
SharedReg806_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg806_out;
SharedReg930_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg930_out;
SharedReg805_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg805_out;
SharedReg164_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg164_out;
SharedReg871_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg871_out;
SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg828_out;
SharedReg731_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg731_out;
SharedReg830_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg830_out;
SharedReg831_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg831_out;
   MUX_Product28_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg832_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg736_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg887_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg849_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg883_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg924_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg803_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg896_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg806_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg930_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg805_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg164_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg871_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg828_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg731_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg830_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg831_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg938_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg609_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg729_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg934_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg610_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg915_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg615_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_4_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_0_out,
                 Y => Delay1No152_out);

SharedReg244_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg64_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg64_out;
SharedReg108_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg108_out;
SharedReg425_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg425_out;
SharedReg911_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
SharedReg819_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg819_out;
SharedReg914_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg914_out;
SharedReg730_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg730_out;
SharedReg885_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg886_out;
SharedReg427_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg427_out;
SharedReg117_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg117_out;
SharedReg867_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg867_out;
SharedReg729_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg729_out;
SharedReg928_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg928_out;
SharedReg804_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg804_out;
SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg895_out;
SharedReg421_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg421_out;
SharedReg872_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg872_out;
SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg424_out;
SharedReg909_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg909_out;
SharedReg884_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg884_out;
SharedReg65_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg65_out;
SharedReg241_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg241_out;
SharedReg937_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg937_out;
SharedReg612_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg612_out;
SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg424_out;
   MUX_Product28_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg64_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg886_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg427_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg117_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg867_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg729_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg928_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg804_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg421_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg872_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg108_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg909_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg884_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg65_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg241_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg937_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg612_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg424_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg425_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg911_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg819_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg914_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg730_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg885_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_4_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product213_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_0_impl_out,
                 X => Delay1No154_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast);

SharedReg895_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg895_out;
SharedReg892_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg892_out;
SharedReg872_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg872_out;
SharedReg925_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg925_out;
SharedReg901_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg901_out;
SharedReg884_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg884_out;
SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg72_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg72_out;
SharedReg860_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg860_out;
SharedReg190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg190_out;
SharedReg34_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg34_out;
SharedReg863_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg863_out;
SharedReg130_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg130_out;
SharedReg865_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg865_out;
SharedReg936_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg936_out;
SharedReg911_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg912_out;
SharedReg904_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg904_out;
SharedReg768_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg768_out;
SharedReg906_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg906_out;
SharedReg854_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg854_out;
SharedReg855_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg856_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg856_out;
SharedReg83_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg83_out;
SharedReg867_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg867_out;
SharedReg852_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg852_out;
SharedReg928_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg928_out;
SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg567_out;
   MUX_Product213_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg895_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg892_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg34_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg863_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg130_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg865_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg936_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg911_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg912_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg904_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg768_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg906_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg872_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg854_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg856_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg83_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg867_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg852_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg928_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg925_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg901_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg884_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg72_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg860_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_0_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_0_out,
                 Y => Delay1No154_out);

SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg373_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg373_out;
SharedReg702_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg376_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg376_out;
SharedReg769_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg769_out;
SharedReg73_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg73_out;
SharedReg858_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg859_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg859_out;
SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg861_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg861_out;
SharedReg862_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg862_out;
SharedReg130_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg130_out;
SharedReg864_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg864_out;
SharedReg191_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg191_out;
SharedReg377_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg377_out;
SharedReg372_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg372_out;
SharedReg567_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg567_out;
SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg569_out;
SharedReg914_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg914_out;
SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg569_out;
SharedReg573_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg573_out;
SharedReg706_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg706_out;
SharedReg379_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg379_out;
SharedReg878_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg878_out;
SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg699_out;
SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg699_out;
SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg699_out;
SharedReg929_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg929_out;
   MUX_Product213_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg373_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg862_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg130_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg864_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg191_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg377_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg372_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg567_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg914_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg569_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg702_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg573_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg706_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg379_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg878_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg699_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg929_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg376_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg769_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg73_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg859_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg861_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_0_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product213_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_4_impl_out,
                 X => Delay1No156_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast);

SharedReg66_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg262_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg262_out;
SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg623_out;
SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg623_out;
SharedReg925_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg925_out;
SharedReg860_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg860_out;
SharedReg867_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg867_out;
SharedReg872_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg872_out;
SharedReg895_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg895_out;
SharedReg928_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg928_out;
SharedReg863_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg863_out;
SharedReg901_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg901_out;
SharedReg884_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg884_out;
SharedReg906_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg906_out;
SharedReg865_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg865_out;
SharedReg852_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg852_out;
SharedReg904_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg904_out;
SharedReg911_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg911_out;
SharedReg854_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg854_out;
SharedReg912_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg912_out;
SharedReg856_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg856_out;
SharedReg855_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg855_out;
SharedReg936_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg936_out;
   MUX_Product213_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg262_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg863_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg901_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg884_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg906_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg865_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg852_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg904_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg911_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg854_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg912_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg856_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg855_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg936_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg623_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg925_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg860_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg867_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg872_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg895_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg928_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product213_4_impl_0_LUT_out,
                 oMux => MUX_Product213_4_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_4_impl_0_out,
                 Y => Delay1No156_out);

SharedReg117_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg65_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
SharedReg178_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg178_out;
SharedReg263_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg263_out;
SharedReg817_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg817_out;
SharedReg441_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg441_out;
SharedReg440_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg440_out;
SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg739_out;
SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg739_out;
SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg739_out;
SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg625_out;
SharedReg629_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg629_out;
SharedReg436_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg436_out;
SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg625_out;
SharedReg443_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg443_out;
SharedReg746_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg746_out;
SharedReg623_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg623_out;
SharedReg742_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg742_out;
SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg739_out;
SharedReg929_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg929_out;
SharedReg862_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg862_out;
SharedReg861_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg861_out;
SharedReg858_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg858_out;
   MUX_Product213_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg629_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg436_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg625_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg443_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg746_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg623_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg742_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg929_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg178_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg862_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg861_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg858_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg263_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg817_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg441_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg440_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg739_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product213_4_impl_1_LUT_out,
                 oMux => MUX_Product213_4_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_4_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Subtract16_0_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Subtract16_0_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Subtract16_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_0_impl_out,
                 X => Delay1No158_out_to_Subtract16_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Subtract16_0_impl_parent_implementedSystem_port_1_cast);

SharedReg573_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg573_out;
SharedReg3_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg8_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg280_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg280_out;
SharedReg504_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg504_out;
SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg685_out;
SharedReg198_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg198_out;
SharedReg572_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg572_out;
SharedReg705_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg705_out;
SharedReg72_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg72_out;
SharedReg769_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg769_out;
SharedReg375_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg375_out;
SharedReg458_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg458_out;
SharedReg512_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg512_out;
SharedReg197_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg197_out;
SharedReg538_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg538_out;
SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg685_out;
SharedReg767_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg767_out;
SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg380_out;
SharedReg373_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg373_out;
SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg377_out;
SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg377_out;
SharedReg507_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg507_out;
SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg380_out;
SharedReg277_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg277_out;
SharedReg194_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg194_out;
   MUX_Subtract16_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg573_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg705_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg72_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg769_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg375_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg458_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg512_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg197_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg538_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg767_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg6_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg373_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg377_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg507_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg380_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg277_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg194_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg11_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg280_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg504_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg685_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg198_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg572_out_to_MUX_Subtract16_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_0_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_0_impl_0_out,
                 Y => Delay1No158_out);

SharedReg578_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg578_out;
SharedReg19_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg24_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg507_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg507_out;
SharedReg749_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg749_out;
SharedReg689_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg689_out;
SharedReg132_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg132_out;
SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg580_out;
SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg580_out;
SharedReg187_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg187_out;
SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg699_out;
SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
SharedReg457_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg457_out;
Delay17No25_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_16_cast <= Delay17No25_out;
Delay72No_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_17_cast <= Delay72No_out;
SharedReg688_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg688_out;
SharedReg754_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg754_out;
SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg372_out;
SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg568_out;
SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg372_out;
SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg699_out;
SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg372_out;
SharedReg687_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg687_out;
SharedReg569_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg569_out;
SharedReg454_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg454_out;
SharedReg135_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg135_out;
   MUX_Subtract16_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg578_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg187_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg457_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay17No25_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay72No_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg688_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg754_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg22_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg568_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg699_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg372_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg687_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg569_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg454_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg135_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg27_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg507_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg749_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg689_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg132_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg580_out_to_MUX_Subtract16_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_0_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_0_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Subtract16_1_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Subtract16_1_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Subtract16_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_1_impl_out,
                 X => Delay1No160_out_to_Subtract16_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Subtract16_1_impl_parent_implementedSystem_port_1_cast);

SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg393_out;
SharedReg752_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg396_out;
SharedReg283_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg283_out;
SharedReg212_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg212_out;
SharedReg587_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg587_out;
SharedReg3_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg8_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg286_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg286_out;
SharedReg513_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg513_out;
SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg645_out;
SharedReg216_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg216_out;
SharedReg586_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg586_out;
SharedReg715_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg715_out;
SharedReg83_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg83_out;
SharedReg781_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg781_out;
SharedReg391_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg391_out;
SharedReg468_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg468_out;
SharedReg521_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg521_out;
SharedReg215_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg215_out;
SharedReg545_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg545_out;
SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg645_out;
SharedReg779_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg779_out;
SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg396_out;
SharedReg389_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg389_out;
   MUX_Subtract16_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg393_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg286_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg513_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg216_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg586_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg715_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg83_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg781_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg391_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg752_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg468_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg521_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg215_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg545_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg645_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg779_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg389_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg396_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg283_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg212_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg587_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Subtract16_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_1_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_1_impl_0_out,
                 Y => Delay1No160_out);

SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg709_out;
SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg647_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg647_out;
SharedReg583_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg583_out;
SharedReg464_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg464_out;
SharedReg147_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
SharedReg592_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg592_out;
SharedReg19_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg24_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg516_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg516_out;
SharedReg659_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg659_out;
SharedReg649_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg649_out;
SharedReg144_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg144_out;
SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg594_out;
SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg594_out;
SharedReg205_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg205_out;
SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg709_out;
SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg582_out;
SharedReg467_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg467_out;
Delay17No26_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_22_cast <= Delay17No26_out;
Delay72No1_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_23_cast <= Delay72No1_out;
SharedReg648_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg648_out;
SharedReg664_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg664_out;
SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg388_out;
SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg582_out;
SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg388_out;
   MUX_Subtract16_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg516_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg659_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg649_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg144_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg594_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg205_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg709_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg647_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg467_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay17No26_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay72No1_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg648_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg664_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg582_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg388_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg583_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg464_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg592_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Subtract16_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_1_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_1_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Subtract16_2_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Subtract16_2_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Subtract16_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_2_impl_out,
                 X => Delay1No162_out_to_Subtract16_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Subtract16_2_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg652_out;
SharedReg791_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg791_out;
SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg412_out;
SharedReg405_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg405_out;
SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg409_out;
SharedReg298_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg298_out;
SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg412_out;
SharedReg289_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg289_out;
SharedReg230_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg230_out;
SharedReg601_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg601_out;
SharedReg3_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg11_out;
SharedReg8_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
SharedReg292_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg292_out;
SharedReg295_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg295_out;
SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg652_out;
SharedReg234_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg234_out;
SharedReg600_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg600_out;
SharedReg725_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg725_out;
SharedReg94_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg94_out;
SharedReg793_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg793_out;
SharedReg407_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg407_out;
SharedReg478_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg478_out;
SharedReg303_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg303_out;
SharedReg233_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg233_out;
   MUX_Subtract16_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg230_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg601_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg3_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg11_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg292_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg295_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg652_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg234_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg791_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg600_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg725_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg94_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg793_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg407_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg478_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg303_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg233_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg405_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg409_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg298_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg412_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg289_out_to_MUX_Subtract16_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_2_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_2_impl_0_out,
                 Y => Delay1No162_out);

SharedReg655_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg655_out;
SharedReg673_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg673_out;
SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg596_out;
SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg404_out;
SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg719_out;
SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg404_out;
SharedReg338_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg338_out;
SharedReg597_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg597_out;
SharedReg474_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg474_out;
SharedReg159_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg606_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg606_out;
SharedReg19_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg24_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg24_out;
SharedReg298_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg298_out;
SharedReg668_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg668_out;
SharedReg656_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg656_out;
SharedReg156_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg156_out;
SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg608_out;
SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg608_out;
SharedReg223_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg223_out;
SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg719_out;
SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg596_out;
SharedReg477_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg477_out;
Delay17No27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_27_cast <= Delay17No27_out;
Delay72No2_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_28_cast <= Delay72No2_out;
   MUX_Subtract16_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg655_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg673_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg606_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg24_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg298_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg668_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg656_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg156_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg608_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg223_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg477_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay17No27_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay72No2_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg596_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg719_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg404_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg338_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg597_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg474_out_to_MUX_Subtract16_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_2_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_2_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Subtract16_3_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Subtract16_3_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Subtract16_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_3_impl_out,
                 X => Delay1No164_out_to_Subtract16_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Subtract16_3_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg805_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg805_out;
SharedReg423_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg423_out;
SharedReg488_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg488_out;
SharedReg529_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg529_out;
SharedReg251_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg251_out;
SharedReg552_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg552_out;
SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg637_out;
SharedReg803_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg803_out;
SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg428_out;
SharedReg421_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg421_out;
SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg425_out;
SharedReg671_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg671_out;
SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg428_out;
SharedReg310_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg310_out;
SharedReg248_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg248_out;
SharedReg615_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg615_out;
SharedReg3_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg11_out;
SharedReg8_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg8_out;
SharedReg313_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg313_out;
SharedReg522_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg522_out;
SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg637_out;
SharedReg252_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg252_out;
SharedReg614_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg614_out;
SharedReg735_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg735_out;
   MUX_Subtract16_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg805_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg421_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg425_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg671_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg310_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg248_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg615_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg3_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg6_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg423_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg11_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg8_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg313_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg522_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg252_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg614_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg735_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg488_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg529_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg251_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg552_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg637_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg803_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg428_out_to_MUX_Subtract16_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_3_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_3_impl_0_out,
                 Y => Delay1No164_out);

SharedReg241_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg241_out;
SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg729_out;
SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg610_out;
SharedReg487_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg487_out;
Delay17No28_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_5_cast <= Delay17No28_out;
Delay72No3_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_6_cast <= Delay72No3_out;
SharedReg640_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg640_out;
SharedReg682_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg682_out;
SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg420_out;
SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg610_out;
SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg420_out;
SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg729_out;
SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg420_out;
SharedReg639_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg639_out;
SharedReg611_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg611_out;
SharedReg484_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg484_out;
SharedReg171_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg171_out;
SharedReg620_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg620_out;
SharedReg19_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg27_out;
SharedReg24_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg24_out;
SharedReg525_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg525_out;
SharedReg677_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg677_out;
SharedReg641_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg641_out;
SharedReg168_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg168_out;
SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg622_out;
SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg622_out;
   MUX_Subtract16_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg241_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg729_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg639_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg611_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg484_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg171_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg620_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg19_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg22_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg27_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg24_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg525_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg677_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg641_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg168_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg622_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg487_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay17No28_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay72No3_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg640_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg682_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg420_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg610_out_to_MUX_Subtract16_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_3_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_3_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Subtract16_4_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Subtract16_4_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Subtract16_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_4_impl_out,
                 X => Delay1No166_out_to_Subtract16_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Subtract16_4_impl_parent_implementedSystem_port_1_cast);

SharedReg530_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg530_out;
SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg692_out;
SharedReg270_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg270_out;
SharedReg628_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg628_out;
SharedReg745_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg745_out;
SharedReg116_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg116_out;
SharedReg817_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg817_out;
SharedReg439_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg439_out;
SharedReg499_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg499_out;
SharedReg537_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg537_out;
SharedReg269_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg269_out;
SharedReg560_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg692_out;
SharedReg815_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg815_out;
SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg444_out;
SharedReg437_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg437_out;
SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg441_out;
SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg441_out;
SharedReg532_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg532_out;
SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg444_out;
SharedReg304_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg304_out;
SharedReg266_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg266_out;
SharedReg629_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg629_out;
SharedReg3_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg11_out;
SharedReg8_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg8_out;
SharedReg307_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg307_out;
   MUX_Subtract16_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg530_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg269_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg692_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg815_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg437_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg441_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg532_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg444_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg270_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg304_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg266_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg629_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg3_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg6_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg11_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg8_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg307_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg628_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg745_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg116_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg817_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg439_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg499_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg537_out_to_MUX_Subtract16_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_4_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_4_impl_0_out,
                 Y => Delay1No166_out);

SharedReg758_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg758_out;
SharedReg696_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg696_out;
SharedReg180_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg180_out;
SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg636_out;
SharedReg259_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg259_out;
SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg739_out;
SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg624_out;
SharedReg498_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg498_out;
Delay17No29_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_10_cast <= Delay17No29_out;
Delay72No4_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_11_cast <= Delay72No4_out;
SharedReg695_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg695_out;
SharedReg763_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg763_out;
SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg436_out;
SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg624_out;
SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg436_out;
SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg739_out;
SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg436_out;
SharedReg355_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg355_out;
SharedReg625_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg625_out;
SharedReg495_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg495_out;
SharedReg183_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg183_out;
SharedReg634_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg634_out;
SharedReg19_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg19_out;
SharedReg22_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg27_out;
SharedReg24_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg24_out;
SharedReg532_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg532_out;
   MUX_Subtract16_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg758_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg696_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay72No4_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg695_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg763_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg436_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg355_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg625_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg180_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg495_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg183_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg634_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg19_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg22_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg27_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg24_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg532_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg636_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg259_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg739_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg624_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg498_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay17No29_out_to_MUX_Subtract16_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract16_4_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_4_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product316_0_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product316_0_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product316_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product316_0_impl_out,
                 X => Delay1No168_out_to_Product316_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product316_0_impl_parent_implementedSystem_port_1_cast);

SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg767_out;
SharedReg896_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg896_out;
SharedReg770_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg770_out;
SharedReg930_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg930_out;
SharedReg769_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg769_out;
SharedReg128_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg128_out;
SharedReg935_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg935_out;
SharedReg828_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg828_out;
SharedReg701_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg701_out;
SharedReg830_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg830_out;
SharedReg831_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg831_out;
SharedReg832_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg832_out;
SharedReg833_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg833_out;
SharedReg865_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg865_out;
SharedReg938_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg938_out;
SharedReg567_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg567_out;
SharedReg699_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg699_out;
SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg904_out;
SharedReg568_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg568_out;
SharedReg915_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg915_out;
SharedReg573_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg573_out;
SharedReg706_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg706_out;
SharedReg887_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg887_out;
SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg904_out;
SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg767_out;
SharedReg883_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg883_out;
SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg767_out;
SharedReg924_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg924_out;
   MUX_Product316_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg896_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg831_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg832_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg833_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg865_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg938_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg567_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg699_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg568_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg915_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg770_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg573_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg706_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg887_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg904_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg883_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg767_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg924_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg930_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg769_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg935_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg828_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg701_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg830_out_to_MUX_Product316_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product316_0_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_0_impl_0_out,
                 Y => Delay1No168_out);

SharedReg895_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg895_out;
SharedReg373_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg373_out;
SharedReg872_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg872_out;
SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg376_out;
SharedReg909_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg909_out;
SharedReg884_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg884_out;
SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg699_out;
SharedReg187_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg187_out;
SharedReg937_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg570_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg570_out;
SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg376_out;
SharedReg190_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg190_out;
SharedReg192_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg192_out;
SharedReg75_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg75_out;
SharedReg377_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg377_out;
SharedReg911_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg912_out;
SharedReg568_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg568_out;
SharedReg914_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg914_out;
SharedReg700_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg700_out;
SharedReg885_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg886_out;
SharedReg379_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg379_out;
SharedReg709_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg709_out;
SharedReg867_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg867_out;
SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg699_out;
SharedReg928_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg928_out;
SharedReg768_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg768_out;
   MUX_Product316_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg895_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg373_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg190_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg192_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg75_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg377_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg911_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg912_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg568_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg914_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg700_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg872_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg885_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg886_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg379_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg709_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg867_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg928_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg768_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg376_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg909_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg884_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg699_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg187_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg570_out_to_MUX_Product316_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product316_0_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_0_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product316_4_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product316_4_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product316_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product316_4_impl_out,
                 X => Delay1No170_out_to_Product316_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product316_4_impl_parent_implementedSystem_port_1_cast);

SharedReg176_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg817_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg817_out;
SharedReg741_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg741_out;
SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg815_out;
SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg815_out;
SharedReg629_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg629_out;
SharedReg623_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg623_out;
SharedReg746_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg746_out;
SharedReg739_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg739_out;
SharedReg818_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg818_out;
SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg815_out;
SharedReg930_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg930_out;
SharedReg924_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg924_out;
SharedReg915_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg915_out;
SharedReg883_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg883_out;
SharedReg904_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg904_out;
SharedReg887_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg887_out;
SharedReg865_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg865_out;
SharedReg832_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg832_out;
SharedReg831_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg831_out;
SharedReg830_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg830_out;
SharedReg935_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg935_out;
SharedReg938_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg938_out;
   MUX_Product316_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg817_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg930_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg924_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg915_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg883_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg904_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg887_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg865_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg832_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg831_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg741_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg830_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg935_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg938_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg629_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg623_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg746_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg739_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg818_out_to_MUX_Product316_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product316_4_impl_0_LUT_out,
                 oMux => MUX_Product316_4_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_4_impl_0_out,
                 Y => Delay1No170_out);

SharedReg119_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg119_out;
SharedReg262_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg262_out;
SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg440_out;
SharedReg626_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg626_out;
SharedReg441_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg441_out;
SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg739_out;
SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg440_out;
SharedReg816_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg816_out;
SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg739_out;
SharedReg740_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg740_out;
SharedReg443_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg443_out;
SharedReg624_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg624_out;
SharedReg867_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg867_out;
SharedReg872_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg872_out;
SharedReg895_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg895_out;
SharedReg928_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg928_out;
SharedReg909_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg909_out;
SharedReg884_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg884_out;
SharedReg911_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg911_out;
SharedReg885_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg885_out;
SharedReg912_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg912_out;
SharedReg886_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg886_out;
SharedReg937_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg937_out;
   MUX_Product316_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg119_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg262_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg443_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg624_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg867_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg872_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg895_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg928_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg909_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg884_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg911_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg885_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg912_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg886_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg937_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_3 => SharedReg626_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg441_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg440_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg816_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg739_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg740_out_to_MUX_Product316_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product316_4_impl_1_LUT_out,
                 oMux => MUX_Product316_4_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_4_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Subtract22_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_0_impl_out,
                 X => Delay1No172_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg12_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg505_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg505_out;
SharedReg542_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg542_out;
SharedReg576_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg576_out;
SharedReg377_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg377_out;
SharedReg76_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg76_out;
SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg133_out;
SharedReg774_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg774_out;
SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg189_out;
SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg195_out;
SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg749_out;
SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg749_out;
SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg131_out;
Delay45No_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast <= Delay45No_out;
SharedReg777_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg777_out;
SharedReg188_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg188_out;
SharedReg707_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg707_out;
SharedReg73_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg73_out;
SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg131_out;
SharedReg32_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg32_out;
SharedReg539_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg539_out;
SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg133_out;
SharedReg685_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg685_out;
SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg195_out;
   MUX_Subtract22_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg774_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg749_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay45No_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg777_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg188_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg13_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg707_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg73_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg131_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg32_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg539_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg133_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg685_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg505_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg542_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg576_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg377_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg76_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_0_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_0_impl_0_out,
                 Y => Delay1No172_out);

SharedReg39_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg30_out;
SharedReg28_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg750_out;
SharedReg753_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg753_out;
SharedReg378_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg378_out;
SharedReg387_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg387_out;
SharedReg199_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg199_out;
SharedReg138_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg138_out;
SharedReg580_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg580_out;
SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg187_out;
SharedReg203_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg203_out;
SharedReg689_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg689_out;
SharedReg687_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg687_out;
SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg187_out;
SharedReg461_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg461_out;
Delay74No_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast <= Delay74No_out;
SharedReg32_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg32_out;
SharedReg700_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg700_out;
SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg127_out;
SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg127_out;
SharedReg188_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg188_out;
SharedReg751_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg751_out;
SharedReg74_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg74_out;
SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg750_out;
SharedReg130_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg130_out;
   MUX_Subtract22_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg138_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg580_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg203_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg689_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg687_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg187_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg461_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay74No_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg32_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg29_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg700_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg127_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg188_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg751_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg74_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg130_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg750_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg753_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg378_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg387_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg199_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_0_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_0_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Subtract22_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_1_impl_out,
                 X => Delay1No174_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast);

SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg40_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg546_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg546_out;
SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg645_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg645_out;
SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg213_out;
SharedReg146_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg146_out;
SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg14_out;
SharedReg12_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg514_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg514_out;
SharedReg549_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg549_out;
SharedReg590_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg590_out;
SharedReg393_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg393_out;
SharedReg87_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg87_out;
SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg145_out;
SharedReg786_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg786_out;
SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg207_out;
SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg213_out;
SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg659_out;
SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg659_out;
SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg143_out;
Delay45No1_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast <= Delay45No1_out;
SharedReg789_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg789_out;
SharedReg206_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg206_out;
SharedReg717_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg717_out;
SharedReg84_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg84_out;
   MUX_Subtract22_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg514_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg549_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg590_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg393_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg87_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg786_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg546_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg659_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg143_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay45No1_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg789_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg206_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg717_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg84_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg145_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg645_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg213_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg146_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_1_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_1_impl_0_out,
                 Y => Delay1No174_out);

SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg139_out;
SharedReg206_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg206_out;
SharedReg661_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg661_out;
SharedReg85_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg85_out;
SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg660_out;
SharedReg142_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg142_out;
SharedReg47_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg47_out;
SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg30_out;
SharedReg28_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg660_out;
SharedReg663_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg663_out;
SharedReg394_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg394_out;
SharedReg403_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg403_out;
SharedReg217_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg217_out;
SharedReg150_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg150_out;
SharedReg594_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg594_out;
SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg205_out;
SharedReg221_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg221_out;
SharedReg649_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg649_out;
SharedReg647_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg647_out;
SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg205_out;
SharedReg471_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg471_out;
Delay74No1_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast <= Delay74No1_out;
SharedReg40_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg40_out;
SharedReg710_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg710_out;
SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg139_out;
   MUX_Subtract22_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg663_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg394_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg403_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg217_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg150_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg594_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg221_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg661_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg649_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg647_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg205_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg471_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay74No1_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg40_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg710_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg139_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg85_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg660_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg142_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg47_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_1_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_1_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Subtract22_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_2_impl_out,
                 X => Delay1No176_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast);

Delay45No2_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast <= Delay45No2_out;
SharedReg801_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg801_out;
SharedReg224_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg224_out;
SharedReg727_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg727_out;
SharedReg95_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg155_out;
SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg48_out;
SharedReg347_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg347_out;
SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg157_out;
SharedReg652_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg652_out;
SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg231_out;
SharedReg158_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg158_out;
SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg14_out;
SharedReg12_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg12_out;
SharedReg296_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg296_out;
SharedReg350_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg350_out;
SharedReg604_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg604_out;
SharedReg409_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg409_out;
SharedReg98_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg98_out;
SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg157_out;
SharedReg798_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg798_out;
SharedReg225_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg225_out;
SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg231_out;
SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg668_out;
SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg668_out;
SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg155_out;
   MUX_Subtract22_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay45No2_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg801_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg158_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg13_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg12_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg296_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg350_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg604_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg409_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg224_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg98_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg798_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg225_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg231_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg668_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg727_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg95_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg155_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg347_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg157_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg652_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_2_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_2_impl_0_out,
                 Y => Delay1No176_out);

SharedReg481_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg481_out;
Delay74No2_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast <= Delay74No2_out;
SharedReg48_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg720_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg720_out;
SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg151_out;
SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg151_out;
SharedReg224_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg224_out;
SharedReg474_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg474_out;
SharedReg96_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg96_out;
SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg669_out;
SharedReg154_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg154_out;
SharedReg55_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg55_out;
SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg30_out;
SharedReg28_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg28_out;
SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg669_out;
SharedReg672_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg672_out;
SharedReg410_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg410_out;
SharedReg419_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg419_out;
SharedReg235_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg235_out;
SharedReg162_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg162_out;
SharedReg608_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg608_out;
SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg223_out;
SharedReg239_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg239_out;
SharedReg656_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg656_out;
SharedReg654_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg654_out;
SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg223_out;
   MUX_Subtract22_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg481_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay74No2_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg154_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg55_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg29_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg28_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg672_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg410_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg419_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg48_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg235_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg162_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg608_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg239_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg656_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg654_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg720_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg151_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg224_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg474_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg96_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg669_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_2_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_2_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Subtract22_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_3_impl_out,
                 X => Delay1No178_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast);

SharedReg810_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg810_out;
SharedReg243_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg243_out;
SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg249_out;
SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg677_out;
SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg677_out;
SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg167_out;
Delay45No3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast <= Delay45No3_out;
SharedReg813_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg813_out;
SharedReg242_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg242_out;
SharedReg737_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg737_out;
SharedReg106_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg106_out;
SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg167_out;
SharedReg56_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg56_out;
SharedReg553_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg169_out;
SharedReg637_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg637_out;
SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg249_out;
SharedReg170_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg170_out;
SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg14_out;
SharedReg12_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg12_out;
SharedReg523_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg523_out;
SharedReg556_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg556_out;
SharedReg618_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg618_out;
SharedReg425_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg425_out;
SharedReg109_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg109_out;
SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg169_out;
   MUX_Subtract22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg810_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg106_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg56_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg637_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg170_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg13_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg249_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg12_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg523_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg556_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg618_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg425_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg109_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg169_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg677_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg167_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay45No3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg813_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg242_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg737_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_3_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_3_impl_0_out,
                 Y => Delay1No178_out);

SharedReg622_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg622_out;
SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg241_out;
SharedReg257_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg257_out;
SharedReg366_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg366_out;
SharedReg639_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg639_out;
SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg241_out;
SharedReg492_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg492_out;
Delay74No3_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast <= Delay74No3_out;
SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg56_out;
SharedReg730_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg730_out;
SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg163_out;
SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg163_out;
SharedReg242_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg242_out;
SharedReg679_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg679_out;
SharedReg107_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg107_out;
SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg678_out;
SharedReg166_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg166_out;
SharedReg63_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg63_out;
SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg30_out;
SharedReg28_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg28_out;
SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg678_out;
SharedReg681_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg681_out;
SharedReg426_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg426_out;
SharedReg435_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg435_out;
SharedReg253_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg253_out;
SharedReg174_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg174_out;
   MUX_Subtract22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg622_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg163_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg242_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg679_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg107_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg166_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg63_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg29_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg257_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg28_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg678_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg681_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg426_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg435_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg253_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg174_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg366_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg639_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg241_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg492_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay74No3_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg730_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_3_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_3_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Subtract22_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_4_impl_out,
                 X => Delay1No180_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg564_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg564_out;
SharedReg632_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg632_out;
SharedReg441_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg441_out;
SharedReg120_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg120_out;
SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg181_out;
SharedReg822_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg822_out;
SharedReg261_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg267_out;
SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg758_out;
SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg758_out;
SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg179_out;
Delay45No4_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast <= Delay45No4_out;
SharedReg825_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg825_out;
SharedReg260_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg260_out;
SharedReg747_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg747_out;
SharedReg117_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg117_out;
SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg179_out;
SharedReg64_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg64_out;
SharedReg561_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg561_out;
SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg181_out;
SharedReg692_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg692_out;
SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg267_out;
SharedReg182_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg182_out;
SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg15_out;
SharedReg13_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg14_out;
SharedReg12_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg12_out;
SharedReg531_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg531_out;
   MUX_Subtract22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg564_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg632_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay45No4_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg825_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg260_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg747_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg179_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg64_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg561_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg441_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg692_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg182_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg13_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg12_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg531_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg120_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg181_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg822_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg267_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg758_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_4_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_4_impl_0_out,
                 Y => Delay1No180_out);

SharedReg762_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg762_out;
SharedReg442_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg442_out;
SharedReg451_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg271_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg271_out;
SharedReg186_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg636_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg636_out;
SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg259_out;
SharedReg275_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg275_out;
SharedReg696_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg696_out;
SharedReg694_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg694_out;
SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg259_out;
SharedReg503_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg503_out;
Delay74No4_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast <= Delay74No4_out;
SharedReg64_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg64_out;
SharedReg740_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg740_out;
SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg175_out;
SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg175_out;
SharedReg260_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg260_out;
SharedReg495_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg495_out;
SharedReg118_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg118_out;
SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg759_out;
SharedReg178_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg178_out;
SharedReg71_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg71_out;
SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg31_out;
SharedReg29_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg30_out;
SharedReg28_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg28_out;
SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg759_out;
   MUX_Subtract22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg762_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg442_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg503_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay74No4_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg64_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg740_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg175_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg260_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg495_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg118_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg451_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg178_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg71_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg29_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg28_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg759_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg271_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg186_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg636_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg259_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg275_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg696_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg694_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_4_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_4_impl_1_out,
                 Y => Delay1No181_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay19No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay19No_out);

   Delay19No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => Delay19No1_out);

   Delay19No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => Delay19No2_out);

   Delay19No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay19No3_out);

   Delay19No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => Delay19No4_out);

   Delay18No15_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => Delay18No15_out);

   Delay18No16_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => Delay18No16_out);

   Delay18No17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => Delay18No17_out);

   Delay18No18_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => Delay18No18_out);

   Delay18No19_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => Delay18No19_out);

   Delay17No20_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => Delay17No20_out);

   Delay17No21_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => Delay17No21_out);

   Delay17No22_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => Delay17No22_out);

   Delay17No23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => Delay17No23_out);

   Delay17No24_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => Delay17No24_out);

   Delay17No25_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => Delay17No25_out);

   Delay17No26_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => Delay17No26_out);

   Delay17No27_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => Delay17No27_out);

   Delay17No28_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => Delay17No28_out);

   Delay17No29_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => Delay17No29_out);

   Delay27No10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => Delay27No10_out);

   Delay27No11_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => Delay27No11_out);

   Delay27No12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => Delay27No12_out);

   Delay27No13_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => Delay27No13_out);

   Delay27No14_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => Delay27No14_out);

   Delay45No_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => Delay45No_out);

   Delay45No1_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => Delay45No1_out);

   Delay45No2_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => Delay45No2_out);

   Delay45No3_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => Delay45No3_out);

   Delay45No4_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => Delay45No4_out);

   Delay43No_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => Delay43No_out);

   Delay43No1_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => Delay43No1_out);

   Delay43No2_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => Delay43No2_out);

   Delay43No3_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => Delay43No3_out);

   Delay43No4_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => Delay43No4_out);

   Delay72No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => Delay72No_out);

   Delay72No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => Delay72No1_out);

   Delay72No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => Delay72No2_out);

   Delay72No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => Delay72No3_out);

   Delay72No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => Delay72No4_out);

   Delay74No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => Delay74No_out);

   Delay74No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => Delay74No1_out);

   Delay74No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => Delay74No2_out);

   Delay74No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => Delay74No3_out);

   Delay74No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => Delay74No4_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Product32_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product32_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product32_4_impl_0_LUT_out);

   MUX_Product32_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product32_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product32_4_impl_1_LUT_out);

   MUX_Product6_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product6_4_impl_0_LUT_out);

   MUX_Product6_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product6_4_impl_1_LUT_out);

   MUX_Product213_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product213_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product213_4_impl_0_LUT_out);

   MUX_Product213_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product213_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product213_4_impl_1_LUT_out);

   MUX_Product316_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product316_4_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product316_4_impl_0_LUT_out);

   MUX_Product316_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product316_4_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product316_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_2_impl_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_3_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_4_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_0_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_1_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_2_impl_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_3_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_4_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_3_impl_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_4_impl_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_3_impl_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_0_impl_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_1_impl_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_2_impl_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_3_impl_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_4_impl_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_1_impl_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_3_impl_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_4_impl_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_0_impl_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_2_impl_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_3_impl_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_4_impl_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_4_impl_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_2_impl_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_3_impl_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_2_impl_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_3_impl_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_4_impl_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_0_impl_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_4_impl_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_0_impl_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_1_impl_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_2_impl_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_3_impl_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_4_impl_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product316_0_impl_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product316_4_impl_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_0_impl_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_1_impl_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_2_impl_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_3_impl_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_4_impl_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);
end architecture;

