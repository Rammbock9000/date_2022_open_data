--------------------------------------------------------------------------------
--                         ModuloCounter_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_64_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 63 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_9_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid434304_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid434306)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid434304_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid434304_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid434309
--                  (IntAdderAlternative_27_f250_uid434313)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid434309 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid434309 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid434316
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid434316 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid434316 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid434319
--                   (IntAdderClassical_34_f250_uid434321)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid434319 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid434319 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid434304
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid434304 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid434304 is
   component FPAdd_8_23_uid434304_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid434309 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid434316 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid434319 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid434304_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid434309  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid434316  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid434319  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid434304 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid434304  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_64_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iS_61 : in std_logic_vector(33 downto 0);
          iS_62 : in std_logic_vector(33 downto 0);
          iS_63 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
         iS_61 when "111101",
         iS_62 when "111110",
         iS_63 when "111111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_61_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_61_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_61_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_51_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_51_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_51_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid434833
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid434833 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid434833 is
signal XX_m434834 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m434834 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m434834 <= X ;
   YY_m434834 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid434837
--                   (IntAdderClassical_33_f500_uid434839)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid434837 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid434837 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid434833 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid434837 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid434833  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid434837  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid435228_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid435230)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid435228_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid435228_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid435233
--                  (IntAdderAlternative_27_f250_uid435237)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid435233 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid435233 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid435240
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid435240 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid435240 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid435243
--                   (IntAdderClassical_34_f250_uid435245)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid435243 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid435243 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid435228
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid435228 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid435228 is
   component FPAdd_8_23_uid435228_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid435233 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid435240 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid435243 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid435228_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid435233  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid435240  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid435243  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid435228 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid435228  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_48_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_48_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_48_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0110" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0111" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "1000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0011" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0100" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0101" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0110" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0111" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "1000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0011" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0100" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0101" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0011" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0100" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0101" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0110" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0111" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "1000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0001" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0010" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0011" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0100" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0101" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0110" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0111" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "1000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0001" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0010" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0011" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0101" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0110" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0111" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "1000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0001" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0010" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0011" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0101" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0110" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0111" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "1000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0001" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0010" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0110" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0111" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "1000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0001" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0010" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0011" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0100" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0101" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0010" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0011" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0100" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0101" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0110" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0111" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "1000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0001" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0110" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0111" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "1000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0001" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0010" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0011" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0100" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0101" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0101" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0110" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0111" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "1000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0001" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0010" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0011" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0100" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0010" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0011" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0100" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0101" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0110" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0111" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "1000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0001" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0010" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0011" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0100" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0101" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0110" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0111" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "1000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0001" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0011" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0100" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0101" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0110" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0111" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "1000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0001" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0010" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0010" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0011" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0100" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0101" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0110" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0111" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "1000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0001" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0110" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0111" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "1000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0001" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0010" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0011" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0100" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0101" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0110" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0111" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "1000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0001" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0010" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0011" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0100" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0101" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0110" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0111" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "1000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0011" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0100" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0101" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0110" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0111" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "1000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0001" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0010" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0011" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0100" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0101" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0011" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0100" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0101" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0110" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0111" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "1000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0001" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0010" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0010" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0011" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0100" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0101" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0110" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0111" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "1000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0001" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0101" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0110" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0111" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0001" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "1000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0010" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0011" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0100" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0011" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0100" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0101" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0110" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0111" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "1000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0001" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0010" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0110" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0111" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "1000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0001" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0010" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0011" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0100" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0101" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0011" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0100" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0101" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0110" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0111" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "1000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0001" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0010" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0101" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0110" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0111" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "1000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0001" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0010" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0011" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0100" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0101" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0110" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0111" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "1000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0001" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0010" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0011" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0100" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0010" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0011" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0100" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0101" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0110" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0111" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "1000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0001" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0010" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0011" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0100" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0101" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0110" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0111" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "1000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0001" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0011" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0101" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0110" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0111" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "1000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0001" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0010" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0011" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0100" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0101" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0110" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0111" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "1000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0001" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0010" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0110" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0111" when "001000",
      "0000" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "1000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0001" when "011110",
      "0000" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0010" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0011" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0100" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0101" when "111010",
      "0000" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0000" when "000000",
      "0000" when "000001",
      "0110" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0000" when "000111",
      "0000" when "001000",
      "0111" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "1000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0000" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0001" when "011111",
      "0000" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "0000" when "100101",
      "0010" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0011" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0100" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0000" when "110111",
      "0000" when "111000",
      "0000" when "111001",
      "0000" when "111010",
      "0101" when "111011",
      "0000" when "111100",
      "0000" when "111101",
      "0000" when "111110",
      "0000" when "111111",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000110" when "000000",
      "001010" when "000001",
      "101000" when "000010",
      "010100" when "000011",
      "010110" when "000100",
      "110111" when "000101",
      "100100" when "000110",
      "011001" when "000111",
      "011011" when "001000",
      "011100" when "001001",
      "110101" when "001010",
      "111000" when "001011",
      "010001" when "001100",
      "110100" when "001101",
      "010010" when "001110",
      "100101" when "001111",
      "101100" when "010000",
      "011110" when "010001",
      "001110" when "010010",
      "101001" when "010011",
      "000000" when "010100",
      "111001" when "010101",
      "101111" when "010110",
      "001111" when "010111",
      "111100" when "011000",
      "111011" when "011001",
      "100010" when "011010",
      "000000" when "011011",
      "100011" when "011100",
      "100110" when "011101",
      "011000" when "011110",
      "010000" when "011111",
      "110001" when "100000",
      "100111" when "100001",
      "000000" when "100010",
      "101010" when "100011",
      "001101" when "100100",
      "101011" when "100101",
      "110010" when "100110",
      "110000" when "100111",
      "010111" when "101000",
      "110011" when "101001",
      "011010" when "101010",
      "100001" when "101011",
      "010101" when "101100",
      "100000" when "101101",
      "011111" when "101110",
      "101101" when "101111",
      "011101" when "110000",
      "111010" when "110001",
      "000001" when "110010",
      "000011" when "110011",
      "001100" when "110100",
      "001011" when "110101",
      "000111" when "110110",
      "101110" when "110111",
      "110110" when "111000",
      "010011" when "111001",
      "000000" when "111010",
      "000010" when "111011",
      "000101" when "111100",
      "000100" when "111101",
      "001000" when "111110",
      "001001" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000110" when "000000",
      "001010" when "000001",
      "100110" when "000010",
      "011100" when "000011",
      "011000" when "000100",
      "110101" when "000101",
      "100011" when "000110",
      "010110" when "000111",
      "100001" when "001000",
      "100010" when "001001",
      "110010" when "001010",
      "111001" when "001011",
      "010100" when "001100",
      "110110" when "001101",
      "011001" when "001110",
      "100101" when "001111",
      "101110" when "010000",
      "011101" when "010001",
      "001110" when "010010",
      "101000" when "010011",
      "000000" when "010100",
      "001111" when "010101",
      "101101" when "010110",
      "001101" when "010111",
      "010001" when "011000",
      "010000" when "011001",
      "111100" when "011010",
      "000000" when "011011",
      "110111" when "011100",
      "100100" when "011101",
      "111010" when "011110",
      "010011" when "011111",
      "101111" when "100000",
      "100111" when "100001",
      "000000" when "100010",
      "101001" when "100011",
      "010010" when "100100",
      "101010" when "100101",
      "110001" when "100110",
      "110000" when "100111",
      "111011" when "101000",
      "110011" when "101001",
      "010111" when "101010",
      "011110" when "101011",
      "010101" when "101100",
      "100000" when "101101",
      "011111" when "101110",
      "101011" when "101111",
      "011011" when "110000",
      "111000" when "110001",
      "000010" when "110010",
      "000100" when "110011",
      "001100" when "110100",
      "001011" when "110101",
      "000111" when "110110",
      "101100" when "110111",
      "110100" when "111000",
      "011010" when "111001",
      "000001" when "111010",
      "000011" when "111011",
      "000000" when "111100",
      "000101" when "111101",
      "001000" when "111110",
      "001001" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000100" when "000000",
      "000010" when "000001",
      "101011" when "000010",
      "010101" when "000011",
      "001111" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "101001" when "000111",
      "110000" when "001000",
      "001001" when "001001",
      "000111" when "001010",
      "110001" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "011001" when "001110",
      "100000" when "001111",
      "001011" when "010000",
      "101000" when "010001",
      "100011" when "010010",
      "101111" when "010011",
      "000000" when "010100",
      "011111" when "010101",
      "101101" when "010110",
      "001010" when "010111",
      "100110" when "011000",
      "101110" when "011001",
      "001000" when "011010",
      "000000" when "011011",
      "000110" when "011100",
      "100100" when "011101",
      "110010" when "011110",
      "100101" when "011111",
      "101010" when "100000",
      "100010" when "100001",
      "000000" when "100010",
      "010110" when "100011",
      "100111" when "100100",
      "001110" when "100101",
      "011011" when "100110",
      "010100" when "100111",
      "100001" when "101000",
      "000000" when "101001",
      "011000" when "101010",
      "001101" when "101011",
      "001100" when "101100",
      "010011" when "101101",
      "010001" when "101110",
      "010111" when "101111",
      "000000" when "110000",
      "011110" when "110001",
      "010010" when "110010",
      "011101" when "110011",
      "010000" when "110100",
      "011100" when "110101",
      "011010" when "110110",
      "000000" when "110111",
      "000000" when "111000",
      "101100" when "111001",
      "000000" when "111010",
      "000001" when "111011",
      "000101" when "111100",
      "000011" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000100" when "000000",
      "000010" when "000001",
      "101100" when "000010",
      "010011" when "000011",
      "001110" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "101001" when "000111",
      "110010" when "001000",
      "001000" when "001001",
      "000111" when "001010",
      "110001" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "010111" when "001110",
      "100000" when "001111",
      "000110" when "010000",
      "100100" when "010001",
      "100001" when "010010",
      "101111" when "010011",
      "000000" when "010100",
      "011100" when "010101",
      "101110" when "010110",
      "001010" when "010111",
      "100101" when "011000",
      "110000" when "011001",
      "101000" when "011010",
      "000000" when "011011",
      "100111" when "011100",
      "101010" when "011101",
      "001001" when "011110",
      "100011" when "011111",
      "101011" when "100000",
      "100010" when "100001",
      "000000" when "100010",
      "010100" when "100011",
      "100110" when "100100",
      "001100" when "100101",
      "010110" when "100110",
      "010001" when "100111",
      "011111" when "101000",
      "000000" when "101001",
      "010101" when "101010",
      "001011" when "101011",
      "010000" when "101100",
      "011110" when "101101",
      "010010" when "101110",
      "011101" when "101111",
      "000000" when "110000",
      "011010" when "110001",
      "001111" when "110010",
      "011000" when "110011",
      "001101" when "110100",
      "011011" when "110101",
      "011001" when "110110",
      "000000" when "110111",
      "000000" when "111000",
      "101101" when "111001",
      "000000" when "111010",
      "000001" when "111011",
      "000101" when "111100",
      "000011" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000100" when "000000",
      "000011" when "000001",
      "011010" when "000010",
      "001100" when "000011",
      "001101" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "011101" when "000111",
      "010010" when "001000",
      "010011" when "001001",
      "100111" when "001010",
      "101000" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "011001" when "001110",
      "011100" when "001111",
      "101100" when "010000",
      "100011" when "010001",
      "010110" when "010010",
      "000000" when "010011",
      "000000" when "010100",
      "100101" when "010101",
      "101001" when "010110",
      "001000" when "010111",
      "101111" when "011000",
      "101110" when "011001",
      "000000" when "011010",
      "000000" when "011011",
      "000110" when "011100",
      "100001" when "011101",
      "101101" when "011110",
      "101011" when "011111",
      "011111" when "100000",
      "000000" when "100001",
      "000000" when "100010",
      "100000" when "100011",
      "000111" when "100100",
      "100100" when "100101",
      "100010" when "100110",
      "100110" when "100111",
      "011110" when "101000",
      "000000" when "101001",
      "011000" when "101010",
      "001001" when "101011",
      "001010" when "101100",
      "010001" when "101101",
      "001111" when "101110",
      "010100" when "101111",
      "000000" when "110000",
      "010101" when "110001",
      "010000" when "110010",
      "011011" when "110011",
      "001110" when "110100",
      "010111" when "110101",
      "001011" when "110110",
      "000000" when "110111",
      "000000" when "111000",
      "101010" when "111001",
      "000000" when "111010",
      "000001" when "111011",
      "000101" when "111100",
      "000010" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000100" when "000000",
      "000011" when "000001",
      "011010" when "000010",
      "010100" when "000011",
      "001110" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "100000" when "000111",
      "011001" when "001000",
      "011100" when "001001",
      "101010" when "001010",
      "101100" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "010111" when "001110",
      "100001" when "001111",
      "101111" when "010000",
      "101000" when "010001",
      "010101" when "010010",
      "000000" when "010011",
      "000000" when "010100",
      "100110" when "010101",
      "000110" when "010110",
      "001011" when "010111",
      "001001" when "011000",
      "001000" when "011001",
      "000000" when "011010",
      "000000" when "011011",
      "101101" when "011100",
      "100111" when "011101",
      "000111" when "011110",
      "101110" when "011111",
      "100010" when "100000",
      "000000" when "100001",
      "000000" when "100010",
      "100011" when "100011",
      "001010" when "100100",
      "100101" when "100101",
      "100100" when "100110",
      "101001" when "100111",
      "011111" when "101000",
      "000000" when "101001",
      "010110" when "101010",
      "001100" when "101011",
      "010000" when "101100",
      "011110" when "101101",
      "010001" when "101110",
      "011101" when "101111",
      "000000" when "110000",
      "010011" when "110001",
      "001111" when "110010",
      "011000" when "110011",
      "001101" when "110100",
      "011011" when "110101",
      "010010" when "110110",
      "000000" when "110111",
      "000000" when "111000",
      "101011" when "111001",
      "000001" when "111010",
      "000010" when "111011",
      "000101" when "111100",
      "000000" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 42 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      Y <= s41;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      Y <= s32;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_64_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_9_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_64_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iS_61 : in std_logic_vector(33 downto 0);
             iS_62 : in std_logic_vector(33 downto 0);
             iS_63 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_61_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_51_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_48_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount641_out : std_logic_vector(5 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add2_8_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add2_8_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add11_8_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add11_8_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract10_8_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract10_8_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1427_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1425_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1402_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1417_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1418_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1364_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1437_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1456_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1445_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1346_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1453_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1451_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1396_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1399_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1320_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No6_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1391_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1320_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1318_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1473_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1466_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1479_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1481_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1461_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1409_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1419_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1356_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1455_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1330_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No3_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1330_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No4_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1344_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1392_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No5_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1398_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1382_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No6_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1474_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1464_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1459_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No8_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1405_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1411_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1412_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1424_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1406_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1415_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1416_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1352_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1358_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1359_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1402_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1367_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1369_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1359_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1362_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1363_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1357_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1406_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1433_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1439_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1440_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1448_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1450_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1434_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1440_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1443_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1444_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1332_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1333_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1438_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1341_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1327_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1333_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1336_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1337_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1331_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1384_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1385_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1389_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1385_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1388_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1389_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1383_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1482_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1588_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1634_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1486_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1487_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1462_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1489_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1630_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1490_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1603_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1604_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1631_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1467_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1524_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1641_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1635_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1528_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1498_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1499_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1500_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1501_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1502_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1591_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1503_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1504_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1593_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1506_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1507_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1509_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1510_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1560_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1511_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1512_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1513_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1514_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1565_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1621_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1517_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1518_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1519_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1520_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1532_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1521_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1522_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1585_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1523_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1648_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1640_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1594_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1601_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1633_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1628_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1470_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1471_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1465_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1566_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1459_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1476_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1406_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1414_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1408_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1420_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1421_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1402_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1366_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1361_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1355_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1357_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1365_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1446_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1447_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1434_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1442_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1438_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1339_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1340_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1327_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1335_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1434_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1331_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1341_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1387_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1389_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1383_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1393_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product31_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product31_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1379_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1394_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product31_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product31_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1483_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1646_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1485_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1595_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1632_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1616_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1492_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1600_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1494_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1496_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1497_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1574_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1615_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1525_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1526_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1527_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1636_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1552_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1554_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1638_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1508_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1639_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1605_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1561_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1562_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1564_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1515_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1531_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1516_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1569_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1570_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1625_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1533_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1583_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1535_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1571_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1613_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1541_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1542_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1617_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1547_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1550_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1551_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1553_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1597_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1555_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1599_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1556_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1463_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1563_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1465_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1475_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1567_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1568_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1459_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1581_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1572_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1586_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1573_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No9_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1402_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1410_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No10_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1364_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1437_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No11_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1445_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No12_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1453_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No40_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No13_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1345_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1392_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1399_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No41_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No14_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1398_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1390_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No24_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1466_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1473_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1423_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1414_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1408_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1421_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1422_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1408_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1420_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1366_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1368_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1361_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1359_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1355_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1367_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1355_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1365_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1447_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1449_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1442_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1440_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1353_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1351_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1446_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1352_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1448_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1436_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1342_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1335_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1333_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1339_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1433_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1341_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1433_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1325_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1341_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1387_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1326_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1328_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1385_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1381_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1377_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1395_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1386_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1393_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1394_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1378_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1394_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product32_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product32_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1650_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1484_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1539_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1589_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1488_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1649_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1647_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1491_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1545_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1602_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1493_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1495_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1548_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1549_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1614_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1629_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1577_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1467_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1529_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1579_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1642_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1596_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1590_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1598_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1592_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1637_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1505_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1463_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1558_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1645_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1619_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1606_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1607_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1530_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1580_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1608_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1609_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1624_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1610_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1611_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1534_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1584_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1626_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1612_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1536_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1477_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1538_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1651_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1540_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1463_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1461_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1543_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1544_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1546_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1575_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1576_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1578_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1643_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1644_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1557_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1559_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1618_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1620_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1475_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1622_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1623_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1462_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1582_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1627_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1476_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1587_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1537_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Subtract3_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Subtract3_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1320_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No17_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1319_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1329_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1322_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1338_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1330_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1323_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1441_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1346_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1324_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1452_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1417_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1419_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1356_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1349_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1413_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1372_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1350_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1371_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1432_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract9_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract9_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1382_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1374_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1373_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1397_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1376_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1375_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No23_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No42_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No15_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1320_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1409_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1408_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No18_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1427_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1403_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1426_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1400_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1347_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1401_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1429_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1330_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1430_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1360_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No20_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1456_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1431_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1454_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Subtract10_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Subtract10_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1474_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1464_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1459_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1480_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount641_instance: ModuloCounter_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount641_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg66_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg368_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg154_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg368_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg290_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg317_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg343_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg368_out;
SharedReg154_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg396_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg235_out;
SharedReg457_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg457_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg343_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg368_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg235_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg290_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg317_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg343_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg396_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg235_out;
SharedReg457_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg457_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg368_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg235_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg36_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg317_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg290_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg317_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg343_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg396_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg235_out;
SharedReg457_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg457_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg368_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg235_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg66_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg396_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg183_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg290_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg317_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg343_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg396_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg235_out;
SharedReg261_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg368_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg235_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg154_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg66_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg368_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg368_out;
SharedReg183_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg368_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg290_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg317_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg343_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg368_out;
SharedReg154_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg396_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg235_out;
SharedReg457_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg457_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg343_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg368_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg235_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg290_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg290_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg290_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg317_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg343_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg368_out;
SharedReg396_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg396_out;
SharedReg183_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg183_out;
SharedReg261_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg368_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg396_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg183_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg290_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg183_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg235_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg235_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg124_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg66_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg396_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg183_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg66_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg95_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg124_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg396_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg183_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg210_out;
SharedReg261_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg853_out;
SharedReg882_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg910_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg940_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg940_out;
SharedReg1321_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg968_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1027_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1057_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1057_out;
SharedReg1086_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg940_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1027_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1057_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg1400_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1321_out;
SharedReg968_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg968_out;
SharedReg998_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1428_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1321_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg968_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg1400_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1347_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1428_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg1400_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1347_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1428_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg1057_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1057_out;
SharedReg1027_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1027_out;
SharedReg853_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg882_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1347_out;
SharedReg910_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg910_out;
SharedReg940_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg940_out;
SharedReg968_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg968_out;
SharedReg1295_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1295_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1057_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1027_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg853_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg882_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1347_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg910_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg940_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg968_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1295_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg1400_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg910_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg1428_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1428_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg1400_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg998_out;
SharedReg1027_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1027_out;
SharedReg1373_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1428_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1321_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg998_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1027_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg940_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg853_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg853_out;
SharedReg1400_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg882_out;
SharedReg910_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg968_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1027_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1057_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1057_out;
SharedReg1086_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg853_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1400_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg882_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1027_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1057_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg1400_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1321_out;
SharedReg968_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg968_out;
SharedReg998_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1428_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1321_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg968_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg853_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg853_out;
SharedReg882_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg910_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg940_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg940_out;
SharedReg1321_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg968_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1027_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1057_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1057_out;
SharedReg1086_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg853_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg940_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1027_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1057_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg853_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg853_out;
SharedReg1400_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg882_out;
SharedReg910_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg940_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg940_out;
SharedReg968_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1027_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1057_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1057_out;
SharedReg1086_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg853_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1400_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg882_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg940_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1027_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1057_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg1400_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1347_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1428_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg1400_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg910_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg1428_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1373_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1086_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1428_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1321_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg1400_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg882_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1347_out;
SharedReg910_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg940_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg940_out;
SharedReg968_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1027_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1057_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1057_out;
SharedReg1457_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg882_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1347_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg940_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1027_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1057_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg1400_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg998_out;
SharedReg1027_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1027_out;
SharedReg1373_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1457_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1457_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1428_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1321_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1027_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1457_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg1400_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1347_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1347_out;
SharedReg1428_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1428_out;
SharedReg1321_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1321_out;
SharedReg998_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg998_out;
SharedReg1027_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1027_out;
SharedReg1373_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1373_out;
SharedReg1295_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1295_out;
SharedReg1086_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1347_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1428_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1321_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg998_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1027_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1373_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1295_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg305_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg487_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg487_out;
SharedReg870_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg870_out;
SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg864_out;
SharedReg691_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg691_out;
SharedReg686_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg686_out;
SharedReg675_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg675_out;
SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg290_out;
SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg854_out;
SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg853_out;
SharedReg1401_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1401_out;
SharedReg490_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg490_out;
SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg54_out;
SharedReg872_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg872_out;
SharedReg1403_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1403_out;
SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg855_out;
SharedReg56_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg56_out;
SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg673_out;
SharedReg1128_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1128_out;
SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg484_out;
SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg295_out;
SharedReg492_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg492_out;
SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg853_out;
SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg864_out;
SharedReg302_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg302_out;
SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg290_out;
SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg863_out;
SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg855_out;
SharedReg503_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg503_out;
SharedReg52_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg52_out;
SharedReg502_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg502_out;
SharedReg678_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg678_out;
SharedReg861_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg861_out;
SharedReg868_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg868_out;
SharedReg1410_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1410_out;
SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg53_out;
SharedReg291_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg291_out;
SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg854_out;
SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg38_out;
SharedReg871_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg871_out;
SharedReg51_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg51_out;
SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg673_out;
SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg484_out;
SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg295_out;
SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg295_out;
SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg860_out;
SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg860_out;
SharedReg1123_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1123_out;
SharedReg1125_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1125_out;
SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg486_out;
SharedReg1118_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1118_out;
SharedReg500_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg500_out;
SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg863_out;
SharedReg301_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg301_out;
SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg486_out;
SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg486_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg870_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg691_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg686_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg675_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1401_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg490_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg872_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1403_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg56_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1128_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg492_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg853_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg864_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg302_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg290_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg855_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg503_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg52_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg502_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg678_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg861_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg868_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1410_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg291_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg854_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg871_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg51_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg673_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg484_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg295_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg860_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1123_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1125_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1118_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg500_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg863_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg301_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg486_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg487_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg677_out;
SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg865_out;
SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg865_out;
SharedReg496_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg496_out;
SharedReg498_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg498_out;
SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1115_out;
SharedReg50_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg50_out;
SharedReg867_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg867_out;
SharedReg880_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg880_out;
SharedReg1427_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1427_out;
SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg673_out;
SharedReg38_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg38_out;
SharedReg856_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg856_out;
SharedReg877_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg877_out;
SharedReg1425_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1425_out;
SharedReg43_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg43_out;
SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1115_out;
SharedReg497_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg497_out;
SharedReg680_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg680_out;
SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg290_out;
SharedReg484_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg484_out;
SharedReg858_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg858_out;
SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg853_out;
SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg292_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg292_out;
SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg853_out;
SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1404_out;
SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg678_out;
SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg290_out;
SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg490_out;
SharedReg676_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg676_out;
SharedReg881_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg881_out;
SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg853_out;
SharedReg879_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg879_out;
SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg36_out;
SharedReg61_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg61_out;
SharedReg875_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg875_out;
SharedReg308_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg308_out;
SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1404_out;
SharedReg315_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg315_out;
SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1115_out;
SharedReg675_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg675_out;
SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg290_out;
SharedReg854_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg854_out;
SharedReg1402_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1402_out;
SharedReg487_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg487_out;
SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1120_out;
SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg677_out;
SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1120_out;
SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg678_out;
SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg853_out;
SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg36_out;
SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg673_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg865_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg496_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg498_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg50_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg867_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg880_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1427_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg38_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg856_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg877_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1425_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg43_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg497_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg680_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg484_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg858_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg292_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg676_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg881_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg879_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg61_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg875_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg308_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1404_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg315_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1115_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg675_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg290_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg854_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1402_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg487_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1120_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg678_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg853_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg673_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg677_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg507_out;
SharedReg1138_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1138_out;
SharedReg521_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg521_out;
SharedReg1410_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1410_out;
SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg76_out;
SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg507_out;
SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg507_out;
SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg79_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg13_out;
SharedReg508_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg508_out;
SharedReg1417_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1417_out;
SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg893_out;
SharedReg711_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg711_out;
SharedReg706_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg706_out;
SharedReg695_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg695_out;
SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg317_out;
SharedReg883_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg883_out;
SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg882_out;
SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1348_out;
SharedReg511_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg511_out;
SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg320_out;
SharedReg1418_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1418_out;
SharedReg1350_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1350_out;
SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg884_out;
SharedReg309_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg309_out;
SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg693_out;
SharedReg1148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1148_out;
SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg505_out;
SharedReg322_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg322_out;
SharedReg513_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg513_out;
SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg882_out;
SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg893_out;
SharedReg329_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg329_out;
SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg317_out;
SharedReg892_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg892_out;
SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg884_out;
SharedReg524_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg524_out;
SharedReg82_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg82_out;
SharedReg523_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg523_out;
SharedReg698_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg698_out;
SharedReg890_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg890_out;
SharedReg897_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg897_out;
SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg505_out;
SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg882_out;
SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg505_out;
SharedReg512_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg512_out;
SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg693_out;
SharedReg321_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg321_out;
SharedReg1438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1438_out;
SharedReg112_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg112_out;
SharedReg96_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg96_out;
SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1348_out;
SharedReg319_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg319_out;
SharedReg928_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg928_out;
SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg110_out;
SharedReg713_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg713_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1138_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg508_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1417_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg711_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg521_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg706_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg695_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg883_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg511_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1418_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1350_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1410_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg309_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1148_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg322_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg513_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg893_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg329_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg892_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg884_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg524_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg82_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg523_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg698_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg890_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg897_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg882_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg505_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg512_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg693_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg321_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg112_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg96_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1348_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg507_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg319_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg928_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg713_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg697_out;
SharedReg1140_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1140_out;
SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg698_out;
SharedReg1400_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1400_out;
SharedReg290_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg290_out;
SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg693_out;
SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg693_out;
SharedReg294_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg294_out;
SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg31_out;
SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg697_out;
SharedReg1413_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1413_out;
SharedReg894_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg894_out;
SharedReg517_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg517_out;
SharedReg519_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg519_out;
SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1135_out;
SharedReg80_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg80_out;
SharedReg896_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg896_out;
SharedReg908_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg908_out;
SharedReg1372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1372_out;
SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg693_out;
Delay80No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast <= Delay80No1_out;
SharedReg885_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg885_out;
SharedReg905_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg905_out;
SharedReg1370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1370_out;
SharedReg73_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg73_out;
SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1135_out;
SharedReg518_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg518_out;
SharedReg700_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg700_out;
SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg317_out;
SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg505_out;
SharedReg887_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg887_out;
SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg882_out;
SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg66_out;
SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg319_out;
SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg882_out;
SharedReg1351_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1351_out;
SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg698_out;
SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg317_out;
SharedReg511_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg511_out;
SharedReg696_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg696_out;
SharedReg909_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg909_out;
SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg882_out;
SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1137_out;
SharedReg903_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg903_out;
SharedReg694_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg694_out;
SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1137_out;
SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg505_out;
SharedReg1142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1142_out;
SharedReg92_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg92_out;
SharedReg937_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg937_out;
SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg317_out;
SharedReg118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg118_out;
SharedReg931_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg931_out;
SharedReg361_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg361_out;
SharedReg914_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg914_out;
SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg366_out;
SharedReg1155_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1155_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1140_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg697_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1413_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg894_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg517_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg519_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg80_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg896_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg908_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay80No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg885_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg905_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1400_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg73_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1135_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg518_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg700_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg887_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg290_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1351_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg698_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg511_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg696_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg909_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg882_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg903_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg694_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg505_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1142_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg92_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg937_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg317_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg931_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg693_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg361_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg914_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1155_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg294_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg141_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg911_out;
SharedReg97_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg97_out;
SharedReg958_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg958_out;
SharedReg139_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg733_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg733_out;
SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg528_out;
SharedReg1158_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1158_out;
SharedReg542_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg542_out;
SharedReg892_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg892_out;
SharedReg328_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg328_out;
SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg528_out;
SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg528_out;
SharedReg332_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg332_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg13_out;
SharedReg529_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg529_out;
SharedReg899_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg899_out;
SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg921_out;
SharedReg731_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg731_out;
SharedReg536_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg536_out;
SharedReg715_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg715_out;
SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg343_out;
SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg911_out;
SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg910_out;
SharedReg1429_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1429_out;
SharedReg532_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg532_out;
SharedReg346_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg346_out;
SharedReg1364_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1364_out;
SharedReg1431_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1431_out;
SharedReg912_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg912_out;
SharedReg86_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg86_out;
SharedReg713_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg713_out;
SharedReg1168_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1168_out;
SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg526_out;
SharedReg348_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg348_out;
SharedReg534_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg534_out;
SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg910_out;
SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg921_out;
SharedReg355_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg355_out;
SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg343_out;
SharedReg920_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg920_out;
SharedReg356_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg356_out;
SharedReg732_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg732_out;
SharedReg1437_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1437_out;
SharedReg718_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg718_out;
SharedReg530_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg530_out;
SharedReg353_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg353_out;
SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg526_out;
SharedReg1430_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1430_out;
SharedReg566_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg566_out;
SharedReg140_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg140_out;
SharedReg565_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg565_out;
SharedReg738_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg738_out;
SharedReg1436_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1436_out;
SharedReg955_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg955_out;
SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg547_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg892_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg328_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg332_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg529_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg899_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg731_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg536_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg715_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg97_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg911_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1429_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg532_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg346_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1364_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1431_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg912_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg86_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg713_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg958_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1168_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg348_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg534_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg355_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg343_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg920_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg356_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg139_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg732_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1437_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg718_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg530_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg353_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg526_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1430_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg566_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg140_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg565_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg733_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg738_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1436_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg955_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg547_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg528_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1158_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg542_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg147_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg961_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg961_out;
SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
SharedReg1432_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1432_out;
SharedReg152_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg152_out;
SharedReg1175_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1175_out;
SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg717_out;
SharedReg1160_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1160_out;
SharedReg718_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg718_out;
SharedReg1347_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1347_out;
SharedReg317_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg317_out;
SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg713_out;
SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg713_out;
SharedReg321_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg321_out;
SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg31_out;
SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg717_out;
SharedReg1360_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1360_out;
SharedReg922_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg922_out;
SharedReg538_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg538_out;
SharedReg723_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg723_out;
SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1155_out;
SharedReg109_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg109_out;
SharedReg924_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg924_out;
SharedReg938_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg938_out;
SharedReg1456_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1456_out;
SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg713_out;
Delay80No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast <= Delay80No2_out;
SharedReg913_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg913_out;
SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg935_out;
SharedReg933_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg933_out;
SharedReg102_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg102_out;
SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1155_out;
SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg539_out;
SharedReg720_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg720_out;
SharedReg343_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg343_out;
SharedReg526_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg526_out;
SharedReg915_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg915_out;
SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg910_out;
SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg95_out;
SharedReg345_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg345_out;
SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg910_out;
SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg96_out;
SharedReg1159_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1159_out;
SharedReg919_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg919_out;
SharedReg1158_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1158_out;
SharedReg1156_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1156_out;
Delay91No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast <= Delay91No2_out;
SharedReg714_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg714_out;
SharedReg1325_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1325_out;
SharedReg738_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg738_out;
SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg124_out;
SharedReg553_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg553_out;
SharedReg736_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg736_out;
SharedReg967_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg967_out;
SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg910_out;
SharedReg1177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1177_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1347_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg317_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg321_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg961_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1360_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg922_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg538_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg723_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg109_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg924_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg938_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1456_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg713_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay80No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg913_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg933_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg102_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1155_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1432_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg720_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg343_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg526_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg915_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg95_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg345_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg96_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg152_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1159_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg919_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1158_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1156_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay91No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg714_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1325_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg738_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg553_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1175_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg736_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg967_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg910_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg717_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1160_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg718_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg587_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg587_out;
SharedReg171_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg171_out;
SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg586_out;
SharedReg758_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg758_out;
SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg948_out;
SharedReg983_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg983_out;
SharedReg568_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg568_out;
SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg172_out;
SharedReg369_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg369_out;
SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg941_out;
SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg126_out;
SharedReg986_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg986_out;
SharedReg384_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg384_out;
SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg753_out;
SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg549_out;
SharedReg1178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1178_out;
SharedReg563_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg563_out;
SharedReg920_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg920_out;
SharedReg354_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg354_out;
SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg549_out;
SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg549_out;
SharedReg358_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg358_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg12_out;
SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg13_out;
SharedReg550_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg550_out;
SharedReg927_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg927_out;
SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg951_out;
SharedReg751_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg751_out;
SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg557_out;
SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg735_out;
SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg368_out;
SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg941_out;
SharedReg940_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg940_out;
SharedReg1322_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1322_out;
SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg553_out;
SharedReg371_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg371_out;
SharedReg1445_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1445_out;
SharedReg1324_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1324_out;
SharedReg942_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg942_out;
SharedReg114_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg114_out;
SharedReg733_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg733_out;
SharedReg1188_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1188_out;
SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg547_out;
SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg735_out;
SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg124_out;
SharedReg1175_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1175_out;
SharedReg1189_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1189_out;
SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg951_out;
SharedReg381_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg381_out;
SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg401_out;
SharedReg576_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg576_out;
SharedReg1321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1321_out;
SharedReg979_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg979_out;
SharedReg408_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg408_out;
SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg368_out;
SharedReg978_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg978_out;
SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg409_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg587_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg986_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg384_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg563_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg920_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg354_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg549_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg358_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg758_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg550_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg927_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg751_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg940_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1322_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg371_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1445_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1324_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg942_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg114_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg733_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1188_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg547_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg983_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg735_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1175_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1189_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg951_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg381_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg576_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg979_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg568_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg408_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg368_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg978_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg172_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg369_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg758_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg758_out;
SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg368_out;
SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg574_out;
SharedReg756_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg756_out;
SharedReg997_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg997_out;
SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg940_out;
SharedReg1197_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1197_out;
SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg124_out;
SharedReg179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg179_out;
SharedReg991_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg991_out;
SharedReg416_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg416_out;
SharedReg1325_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1325_out;
SharedReg394_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg394_out;
SharedReg1195_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1195_out;
SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg737_out;
SharedReg1180_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1180_out;
SharedReg738_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg738_out;
SharedReg1428_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1428_out;
SharedReg343_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg343_out;
SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg733_out;
SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg733_out;
SharedReg347_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg347_out;
SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg30_out;
SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg31_out;
SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg737_out;
SharedReg1441_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1441_out;
SharedReg952_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg952_out;
SharedReg559_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg559_out;
SharedReg743_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg743_out;
SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1175_out;
SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg138_out;
SharedReg954_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg954_out;
SharedReg966_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg966_out;
SharedReg1346_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1346_out;
SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg733_out;
Delay80No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast <= Delay80No3_out;
SharedReg943_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg943_out;
SharedReg1453_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1453_out;
SharedReg1451_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1451_out;
SharedReg131_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg131_out;
SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1175_out;
SharedReg560_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg560_out;
SharedReg740_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg740_out;
SharedReg1179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1179_out;
SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1175_out;
SharedReg374_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg374_out;
SharedReg1192_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1192_out;
SharedReg1177_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1177_out;
SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg940_out;
SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg124_out;
SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg154_out;
SharedReg568_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg568_out;
SharedReg1326_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1326_out;
SharedReg1321_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1321_out;
SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg368_out;
SharedReg156_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg156_out;
SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg940_out;
SharedReg125_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg125_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg758_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg416_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1325_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg394_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1195_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1180_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg738_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1428_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg343_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg347_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg30_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg756_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg737_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1441_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg952_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg559_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg743_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg954_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg966_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1346_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg997_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg733_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => Delay80No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg943_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1453_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1451_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg131_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg560_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg740_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1175_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg374_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1192_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1177_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg568_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1326_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1321_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1197_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg368_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg156_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg940_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg125_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg124_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg179_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg991_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg597_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg597_out;
SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg968_out;
SharedReg1009_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1009_out;
SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg1008_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1008_out;
SharedReg195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg195_out;
SharedReg608_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg608_out;
SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg412_out;
SharedReg607_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg607_out;
SharedReg778_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg778_out;
SharedReg1329_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1329_out;
SharedReg1015_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1015_out;
SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg589_out;
SharedReg413_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg413_out;
SharedReg397_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg397_out;
SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg969_out;
SharedReg156_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg156_out;
SharedReg1017_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1017_out;
SharedReg170_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg170_out;
SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg773_out;
SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg570_out;
SharedReg1198_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1198_out;
SharedReg584_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg584_out;
SharedReg950_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg950_out;
SharedReg379_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg379_out;
SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg570_out;
SharedReg1225_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1225_out;
SharedReg383_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg383_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg12_out;
SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg13_out;
SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg571_out;
SharedReg957_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg957_out;
SharedReg979_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg979_out;
SharedReg771_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg771_out;
SharedReg578_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg578_out;
SharedReg755_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg755_out;
SharedReg396_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg396_out;
SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg969_out;
SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg968_out;
SharedReg999_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg999_out;
SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg574_out;
SharedReg399_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg399_out;
SharedReg959_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg959_out;
SharedReg158_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg158_out;
SharedReg568_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg568_out;
SharedReg401_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg401_out;
SharedReg579_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg579_out;
SharedReg1195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1195_out;
SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg415_out;
SharedReg1018_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1018_out;
SharedReg1030_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1030_out;
SharedReg1000_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1000_out;
SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg174_out;
SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg773_out;
SharedReg1228_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1228_out;
SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg589_out;
SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg589_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg597_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg778_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1329_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1015_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg413_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg397_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg156_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1017_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg170_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1009_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1198_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg584_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg950_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg379_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg570_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1225_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg383_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg957_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg979_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg771_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg578_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg755_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg396_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg969_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg968_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg999_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg399_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg959_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1008_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg158_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg568_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg401_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg579_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1018_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1030_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1000_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg195_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg773_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1228_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg589_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg608_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg607_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg589_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg973_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg973_out;
SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg968_out;
SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg154_out;
SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg398_out;
SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg155_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg778_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg778_out;
SharedReg396_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg396_out;
SharedReg595_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg595_out;
SharedReg776_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg776_out;
SharedReg1056_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1056_out;
SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg968_out;
SharedReg1217_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1217_out;
SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg154_out;
SharedReg206_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg206_out;
SharedReg1050_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1050_out;
SharedReg445_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg445_out;
SharedReg1002_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1002_out;
SharedReg424_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg424_out;
SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1215_out;
SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg757_out;
SharedReg1200_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1200_out;
SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg758_out;
SharedReg1321_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1321_out;
SharedReg368_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg368_out;
SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg753_out;
SharedReg1220_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1220_out;
SharedReg372_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg372_out;
SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg30_out;
SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg31_out;
SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg757_out;
SharedReg1334_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1334_out;
SharedReg980_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg980_out;
SharedReg580_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg580_out;
SharedReg763_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg763_out;
SharedReg1195_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1195_out;
SharedReg169_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg169_out;
SharedReg982_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg982_out;
SharedReg996_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg996_out;
SharedReg1026_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1026_out;
SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg753_out;
Delay80No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast <= Delay80No4_out;
SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1001_out;
SharedReg150_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg150_out;
SharedReg754_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg754_out;
SharedReg392_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg392_out;
SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg585_out;
SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg758_out;
SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg398_out;
SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1001_out;
SharedReg993_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg993_out;
SharedReg1024_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1024_out;
SharedReg190_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg190_out;
SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1215_out;
SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg602_out;
SharedReg780_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg780_out;
SharedReg1219_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1219_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg973_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg776_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1056_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1217_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg206_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1050_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg445_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1002_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg424_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1200_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1321_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg368_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1220_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg372_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg154_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg30_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg757_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1334_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg980_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg580_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg763_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1195_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg169_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg982_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg996_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1026_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg753_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => Delay80No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg968_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg150_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg754_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg392_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg398_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1001_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg993_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1024_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg190_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg155_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1215_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg780_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1219_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg778_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg396_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg595_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_5_impl_out,
                 X => Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1376_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1376_out;
SharedReg1029_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1029_out;
SharedReg417_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg793_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg793_out;
SharedReg1248_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1248_out;
SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg610_out;
SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg610_out;
SharedReg618_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg618_out;
SharedReg1027_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1027_out;
SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1037_out;
SharedReg438_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg438_out;
SharedReg183_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg183_out;
SharedReg1036_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1036_out;
SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg439_out;
SharedReg629_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg629_out;
SharedReg200_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg200_out;
SharedReg628_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg628_out;
SharedReg798_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg798_out;
SharedReg1006_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1006_out;
SharedReg1042_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1042_out;
SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg610_out;
SharedReg201_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg201_out;
SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg427_out;
SharedReg1028_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1028_out;
SharedReg185_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg185_out;
SharedReg1045_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1045_out;
SharedReg199_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg199_out;
SharedReg1066_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1066_out;
SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg591_out;
SharedReg1218_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1218_out;
SharedReg605_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg605_out;
SharedReg978_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg978_out;
SharedReg407_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg407_out;
SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg591_out;
SharedReg1245_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1245_out;
SharedReg411_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg411_out;
SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg12_out;
SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg13_out;
SharedReg592_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg592_out;
SharedReg985_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg985_out;
SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1037_out;
SharedReg791_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg791_out;
SharedReg599_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg599_out;
SharedReg784_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg784_out;
SharedReg1219_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1219_out;
SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg589_out;
SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg589_out;
SharedReg1215_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1215_out;
SharedReg779_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg779_out;
SharedReg806_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg806_out;
SharedReg795_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg795_out;
SharedReg210_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg210_out;
SharedReg1374_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1374_out;
SharedReg1373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1373_out;
SharedReg1058_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1058_out;
SharedReg616_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg616_out;
SharedReg213_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg213_out;
SharedReg1046_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1046_out;
   MUX_Add2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1376_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1029_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg438_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg183_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1036_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg629_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg200_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg628_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg798_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1006_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1042_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg417_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg201_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1028_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg185_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1045_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg199_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1066_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1218_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg793_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg605_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg978_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg407_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg591_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1245_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg411_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg5_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1248_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg7_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg592_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg985_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg791_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg599_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg784_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1219_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg589_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1215_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg779_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg806_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg795_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg210_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1374_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg610_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1058_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg616_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg213_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1046_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg618_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1027_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1037_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_5_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_0_out,
                 Y => Delay1No42_out);

SharedReg1052_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1052_out;
SharedReg1396_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1396_out;
SharedReg433_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg433_out;
SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1235_out;
SharedReg623_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg623_out;
SharedReg800_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg800_out;
SharedReg1239_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1239_out;
SharedReg610_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg610_out;
SharedReg1003_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1003_out;
SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1027_out;
SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg183_out;
SharedReg428_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg428_out;
SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1027_out;
SharedReg184_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg184_out;
SharedReg798_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg798_out;
SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg426_out;
SharedReg616_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg616_out;
SharedReg796_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg796_out;
SharedReg1399_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1399_out;
SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1027_out;
SharedReg1237_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1237_out;
SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg183_out;
SharedReg231_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg231_out;
SharedReg1079_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1079_out;
SharedReg227_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg227_out;
SharedReg1377_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1377_out;
SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg453_out;
SharedReg1083_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1083_out;
SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg777_out;
SharedReg1220_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1220_out;
SharedReg778_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg778_out;
SharedReg998_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg998_out;
SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg154_out;
SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg773_out;
SharedReg1240_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1240_out;
SharedReg400_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg400_out;
SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg30_out;
SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg31_out;
SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg777_out;
SharedReg1011_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1011_out;
SharedReg1039_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1039_out;
SharedReg601_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg601_out;
SharedReg783_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg783_out;
SharedReg1224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1224_out;
SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg773_out;
SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg773_out;
SharedReg596_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg596_out;
SharedReg781_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg781_out;
SharedReg1215_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1215_out;
SharedReg624_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg624_out;
SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1235_out;
SharedReg224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg224_out;
SharedReg1073_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1073_out;
SharedReg1084_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1084_out;
SharedReg1320_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1320_out;
SharedReg793_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg793_out;
Delay80No6_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast <= Delay80No6_out;
SharedReg1376_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1376_out;
   MUX_Add2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1052_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1396_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg428_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg184_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg798_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg616_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg796_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1399_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg433_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1237_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg231_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1079_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg227_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1377_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1083_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1220_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg778_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg998_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1240_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg400_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg23_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg623_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg25_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg30_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg777_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1011_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1039_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg601_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg783_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg800_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg773_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg596_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg781_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1215_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg624_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1235_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg224_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1073_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1084_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1239_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1320_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg793_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => Delay80No6_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1376_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg610_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1003_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1027_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_5_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_6_impl_out,
                 X => Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1058_out;
SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1057_out;
SharedReg1296_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1296_out;
SharedReg637_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg637_out;
SharedReg238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg1076_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1076_out;
SharedReg1060_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1060_out;
SharedReg1059_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1059_out;
SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg446_out;
SharedReg813_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg1268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1268_out;
SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg631_out;
SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg631_out;
SharedReg639_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg639_out;
SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1057_out;
SharedReg1067_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1067_out;
SharedReg247_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg247_out;
SharedReg210_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg210_out;
SharedReg1066_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1066_out;
SharedReg248_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg248_out;
SharedReg650_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg650_out;
SharedReg442_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg442_out;
SharedReg649_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg649_out;
SharedReg818_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg818_out;
SharedReg1381_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1381_out;
SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1074_out;
SharedReg1305_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1305_out;
SharedReg226_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg226_out;
SharedReg236_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg236_out;
SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1058_out;
SharedReg212_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg212_out;
SharedReg1391_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1391_out;
SharedReg225_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg225_out;
SharedReg1102_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1102_out;
SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg612_out;
SharedReg1238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1238_out;
SharedReg626_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg626_out;
SharedReg1036_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1036_out;
SharedReg437_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg437_out;
SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg612_out;
SharedReg1265_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1265_out;
SharedReg441_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg441_out;
SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg8_out;
SharedReg1242_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1242_out;
SharedReg630_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg630_out;
SharedReg220_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg220_out;
SharedReg1254_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1254_out;
SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg13_out;
SharedReg634_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg634_out;
SharedReg1075_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1075_out;
SharedReg1097_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1097_out;
SharedReg831_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg831_out;
SharedReg641_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg641_out;
SharedReg824_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg824_out;
   MUX_Add2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg631_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg639_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1067_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg247_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg210_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1066_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1057_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg248_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg650_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg442_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg649_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg818_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1381_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1305_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg226_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg236_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1296_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1058_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg212_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1391_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg225_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1102_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg626_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1036_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg437_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg637_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg612_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1265_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg441_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg2_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg5_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg238_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1242_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg630_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg220_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1254_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg13_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg634_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1075_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1076_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1097_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg831_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg641_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg824_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1060_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1059_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_6_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_0_out,
                 Y => Delay1No44_out);

SharedReg277_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg1101_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1101_out;
SharedReg1320_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1320_out;
SharedReg1113_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg813_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg813_out;
SharedReg288_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg288_out;
SharedReg1060_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1060_out;
SharedReg1081_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1081_out;
SharedReg1318_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1318_out;
SharedReg217_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg217_out;
SharedReg1255_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1255_out;
SharedReg644_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg644_out;
SharedReg820_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg820_out;
SharedReg1259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1259_out;
SharedReg631_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg631_out;
SharedReg1378_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1378_out;
SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1057_out;
SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg210_out;
SharedReg237_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg237_out;
SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1057_out;
SharedReg211_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg211_out;
SharedReg818_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg818_out;
SharedReg235_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg235_out;
SharedReg637_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg637_out;
SharedReg816_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg816_out;
SharedReg1085_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1085_out;
SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1057_out;
SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1086_out;
SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg210_out;
SharedReg283_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg283_out;
SharedReg1316_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1316_out;
SharedReg254_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg254_out;
SharedReg1299_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1299_out;
SharedReg259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg259_out;
SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1086_out;
SharedReg797_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg797_out;
SharedReg1240_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1240_out;
SharedReg798_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg798_out;
SharedReg1373_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1373_out;
SharedReg183_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg183_out;
SharedReg793_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg793_out;
SharedReg1260_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1260_out;
SharedReg430_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg430_out;
SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg26_out;
SharedReg802_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg802_out;
SharedReg806_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg806_out;
SharedReg222_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg222_out;
SharedReg1248_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1248_out;
SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg31_out;
SharedReg817_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg817_out;
SharedReg1308_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1308_out;
SharedReg1099_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1099_out;
SharedReg643_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg643_out;
SharedReg823_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg823_out;
SharedReg1264_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1264_out;
   MUX_Add2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1101_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1255_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg644_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg820_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg631_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1378_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg237_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1320_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg211_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg818_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg235_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg637_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg816_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1085_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1057_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg210_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg283_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1316_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg254_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1299_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg259_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1086_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg797_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1240_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg798_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1373_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg183_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg813_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg793_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1260_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg430_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg288_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg802_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg806_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg222_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1248_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg31_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg817_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1308_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1060_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1099_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg643_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg823_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1264_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1081_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1318_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg217_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_6_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add2_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_7_impl_out,
                 X => Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1259_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1259_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg631_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg631_out;
SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1255_out;
SharedReg819_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg819_out;
SharedReg851_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg851_out;
SharedReg846_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg846_out;
SharedReg214_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg214_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg631_out;
SharedReg215_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg215_out;
SharedReg642_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg642_out;
SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1255_out;
SharedReg658_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg658_out;
SharedReg474_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg474_out;
SharedReg815_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg815_out;
SharedReg210_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg210_out;
SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1255_out;
SharedReg1269_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1269_out;
SharedReg1067_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1067_out;
SharedReg248_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg248_out;
SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg652_out;
SharedReg832_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg832_out;
SharedReg1304_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1304_out;
SharedReg818_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg818_out;
SharedReg635_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg635_out;
SharedReg245_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg245_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg631_out;
SharedReg469_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg469_out;
SharedReg1057_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1057_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg631_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg631_out;
SharedReg638_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg638_out;
SharedReg813_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg813_out;
SharedReg239_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg239_out;
SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg652_out;
SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg631_out;
SharedReg240_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg240_out;
SharedReg431_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg431_out;
SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1380_out;
SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1380_out;
SharedReg1263_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1263_out;
SharedReg278_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg278_out;
SharedReg1237_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1237_out;
SharedReg1_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg11_out;
SharedReg633_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg633_out;
SharedReg250_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg250_out;
SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg8_out;
SharedReg1262_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1262_out;
SharedReg651_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg651_out;
SharedReg272_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg272_out;
SharedReg1274_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1274_out;
SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg10_out;
   MUX_Add2_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1259_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg642_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg658_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg474_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg815_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg210_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1269_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1067_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg248_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg832_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1304_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg818_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg635_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg245_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg469_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1057_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1255_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg638_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg813_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg239_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg652_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg240_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg431_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1380_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg819_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1263_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg278_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1237_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg3_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg17_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg15_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg11_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg633_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg250_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg851_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg2_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg5_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg16_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg8_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1262_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg651_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg846_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg272_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1274_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg7_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg10_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg214_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg631_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg215_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_7_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_7_impl_0_out,
                 Y => Delay1No46_out);

SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg813_out;
SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg813_out;
SharedReg638_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg638_out;
SharedReg821_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg821_out;
SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1255_out;
SharedReg664_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg664_out;
SharedReg666_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg666_out;
SharedReg233_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg233_out;
SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg814_out;
SharedReg257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg257_out;
SharedReg648_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg648_out;
SharedReg818_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg833_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg833_out;
SharedReg237_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg237_out;
SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1255_out;
SharedReg241_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg241_out;
SharedReg1272_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1272_out;
SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1257_out;
SharedReg1057_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1057_out;
SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg235_out;
SharedReg840_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg840_out;
SharedReg1259_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1259_out;
SharedReg1065_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1065_out;
SharedReg1258_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1258_out;
SharedReg1256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1256_out;
Delay91No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast <= Delay91No7_out;
SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg814_out;
SharedReg457_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg457_out;
SharedReg1108_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1108_out;
SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg814_out;
SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1257_out;
SharedReg631_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg631_out;
SharedReg1262_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1262_out;
SharedReg256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg256_out;
SharedReg834_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg834_out;
SharedReg815_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg815_out;
SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg235_out;
SharedReg1058_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1058_out;
SharedReg1297_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1297_out;
SharedReg634_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg634_out;
SharedReg482_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg482_out;
SharedReg1236_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1236_out;
SharedReg19_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_48_cast <= SharedReg29_out;
SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg813_out;
SharedReg239_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg239_out;
SharedReg18_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_53_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_55_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg26_out;
SharedReg822_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg822_out;
SharedReg826_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_60_cast <= SharedReg826_out;
SharedReg274_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg274_out;
SharedReg1268_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1268_out;
SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg28_out;
   MUX_Add2_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg648_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg833_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg237_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg241_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1272_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1057_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg638_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg840_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1259_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1065_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1258_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay91No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg457_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1108_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg821_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg631_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1262_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg256_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg834_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg815_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg235_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1058_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1297_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1255_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg634_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg482_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1236_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg19_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg21_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg35_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg33_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg29_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg813_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg239_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg664_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg18_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg23_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg30_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg34_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg26_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg822_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg826_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg666_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg274_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1268_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg25_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg233_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg814_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg257_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_7_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_7_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add2_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_8_impl_out,
                 X => Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg1_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg3_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg5_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg11_out;
SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg12_out;
SharedReg13_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg15_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg17_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg251_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg251_out;
SharedReg833_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg833_out;
SharedReg1086_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1086_out;
SharedReg670_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg670_out;
SharedReg839_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg839_out;
SharedReg1473_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1473_out;
SharedReg471_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg471_out;
SharedReg1104_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1104_out;
SharedReg647_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg647_out;
SharedReg1466_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1466_out;
SharedReg1105_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1105_out;
SharedReg279_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg279_out;
SharedReg835_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg835_out;
SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg633_out;
SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg457_out;
SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1087_out;
SharedReg1283_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1283_out;
SharedReg476_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg476_out;
SharedReg246_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg246_out;
SharedReg1066_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1066_out;
SharedReg1258_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1258_out;
SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg457_out;
SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1088_out;
SharedReg662_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg662_out;
SharedReg1460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1460_out;
SharedReg671_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg671_out;
SharedReg1303_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1303_out;
SharedReg655_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg655_out;
SharedReg1288_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1288_out;
SharedReg1096_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1096_out;
SharedReg458_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg458_out;
SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1088_out;
SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg633_out;
SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg654_out;
SharedReg660_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg660_out;
SharedReg263_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg263_out;
SharedReg838_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg838_out;
SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1087_out;
SharedReg460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg460_out;
SharedReg264_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg264_out;
SharedReg1295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1295_out;
SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg654_out;
SharedReg1294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1294_out;
SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1087_out;
SharedReg461_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg461_out;
SharedReg1257_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1257_out;
SharedReg468_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg468_out;
SharedReg1097_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1097_out;
   MUX_Add2_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_61_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg251_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg833_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1086_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg670_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg839_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1473_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg471_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1104_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg647_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1466_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1105_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg279_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg835_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1283_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg3_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg476_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg246_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1066_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1258_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg457_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg662_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg671_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1303_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg655_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1288_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1096_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg458_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1088_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg633_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg660_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg263_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg838_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg5_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg460_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg264_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg654_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1087_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg461_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1257_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg468_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg9_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1097_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_7 => SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_8_impl_0_LUT_out,
                 oMux => MUX_Add2_8_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_8_impl_0_out,
                 Y => Delay1No48_out);

SharedReg23_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg18_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg19_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg21_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg29_out;
SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg30_out;
SharedReg31_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg31_out;
SharedReg33_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg33_out;
SharedReg35_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg35_out;
SharedReg1300_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1300_out;
SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1275_out;
SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg457_out;
SharedReg235_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg235_out;
SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1295_out;
SharedReg261_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg261_out;
SharedReg658_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg658_out;
SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1275_out;
SharedReg818_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg818_out;
SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1275_out;
SharedReg817_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg817_out;
SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1468_out;
SharedReg1298_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1298_out;
SharedReg265_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg265_out;
SharedReg655_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg655_out;
SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1468_out;
SharedReg242_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg242_out;
SharedReg1260_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1260_out;
SharedReg210_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg210_out;
SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1295_out;
SharedReg472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg472_out;
SharedReg1472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1472_out;
SharedReg843_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg843_out;
SharedReg838_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg838_out;
SharedReg1110_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1110_out;
SharedReg837_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg837_out;
SharedReg1114_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1114_out;
SharedReg665_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg665_out;
SharedReg1112_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1112_out;
SharedReg283_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg283_out;
SharedReg813_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg813_out;
SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg833_out;
SharedReg652_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg652_out;
SharedReg1479_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1479_out;
SharedReg836_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg836_out;
SharedReg475_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg475_out;
SharedReg1108_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1108_out;
SharedReg1113_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1113_out;
SharedReg285_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg285_out;
SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg833_out;
SharedReg1288_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1288_out;
Delay80No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_55_cast <= Delay80No8_out;
SharedReg1090_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1090_out;
SharedReg1256_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1256_out;
SharedReg1481_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1481_out;
SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg457_out;
SharedReg1461_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1461_out;
SharedReg459_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg459_out;
   MUX_Add2_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_61_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg31_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg33_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg35_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1300_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg235_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg261_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg658_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg19_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg818_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1275_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg817_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1298_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg265_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg655_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1468_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg242_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1260_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg210_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1295_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1472_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg843_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg838_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1110_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg837_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1114_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg21_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg665_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1112_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg283_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg813_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg652_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1479_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg836_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg475_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1108_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1113_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg285_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg833_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1288_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay80No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1090_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1256_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1481_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg457_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1461_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg27_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg459_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_7 => SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg30_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_8_impl_1_LUT_out,
                 oMux => MUX_Add2_8_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_8_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1117_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1117_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg1122_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1122_out;
SharedReg504_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg504_out;
SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg1134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1134_out;
SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg494_out;
SharedReg684_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg684_out;
SharedReg1119_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1119_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg484_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg484_out;
SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1115_out;
SharedReg679_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg679_out;
SharedReg293_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg293_out;
SharedReg873_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg873_out;
SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg294_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg484_out;
SharedReg295_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg295_out;
SharedReg495_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg495_out;
SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1115_out;
SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg307_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg484_out;
SharedReg675_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg675_out;
SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg36_out;
SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1115_out;
SharedReg1129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1129_out;
SharedReg864_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg864_out;
SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg303_out;
SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg303_out;
SharedReg692_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg692_out;
SharedReg1409_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1409_out;
SharedReg678_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg678_out;
SharedReg488_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg488_out;
SharedReg300_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg300_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg484_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg484_out;
SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg853_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg484_out;
SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg484_out;
SharedReg491_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg491_out;
SharedReg673_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg673_out;
SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg294_out;
SharedReg1357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1357_out;
SharedReg83_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg83_out;
SharedReg318_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg318_out;
SharedReg883_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg883_out;
SharedReg68_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg68_out;
SharedReg900_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg900_out;
SharedReg81_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg81_out;
SharedReg693_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg693_out;
SharedReg505_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg505_out;
SharedReg322_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg322_out;
SharedReg71_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg71_out;
SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1407_out;
SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1407_out;
SharedReg1143_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1143_out;
SharedReg1145_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1145_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1117_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg504_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1134_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg684_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1119_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg679_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg293_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg873_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg295_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg495_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg675_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1115_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg864_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg303_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg692_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1409_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg678_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg488_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg300_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg484_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg491_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg673_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg294_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg83_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg318_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg883_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg68_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg900_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg81_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg693_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg505_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg322_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg71_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1407_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1143_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1145_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1122_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No50_out);

SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1116_out;
SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg682_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg682_out;
SharedReg686_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg686_out;
SharedReg48_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg48_out;
SharedReg1128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1128_out;
SharedReg683_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg683_out;
SharedReg1124_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1124_out;
SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg673_out;
SharedReg491_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg491_out;
SharedReg681_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg681_out;
SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1115_out;
Delay80No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast <= Delay80No_out;
SharedReg1403_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1403_out;
SharedReg64_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg64_out;
SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg674_out;
SharedReg313_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg313_out;
SharedReg501_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg501_out;
SharedReg678_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg678_out;
SharedReg68_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg68_out;
SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1119_out;
SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1115_out;
SharedReg296_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg296_out;
SharedReg1132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1132_out;
SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1117_out;
SharedReg1400_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1400_out;
SharedReg290_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg290_out;
SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg37_out;
SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1119_out;
SharedReg862_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg862_out;
SharedReg1118_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1118_out;
SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1116_out;
Delay91No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast <= Delay91No_out;
SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg674_out;
SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1117_out;
SharedReg875_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg875_out;
SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg674_out;
SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1117_out;
SharedReg484_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg484_out;
SharedReg1122_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1122_out;
SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg63_out;
SharedReg907_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg907_out;
SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg66_out;
SharedReg90_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg90_out;
SharedReg903_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg903_out;
SharedReg335_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg335_out;
SharedReg1351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1351_out;
SharedReg341_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg341_out;
SharedReg1135_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1135_out;
SharedReg695_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg695_out;
SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg66_out;
SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg66_out;
SharedReg1401_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1401_out;
SharedReg884_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg884_out;
SharedReg508_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg508_out;
SharedReg1140_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1140_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg686_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1128_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg683_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1124_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg673_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg491_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg681_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay80No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1403_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg64_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg313_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg501_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg678_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg68_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1115_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg296_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1132_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1400_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg290_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1119_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg862_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1118_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1116_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => Delay91No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg875_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg674_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1117_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg484_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1122_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg907_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg90_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg903_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg335_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg341_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1135_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg695_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg66_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1401_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg884_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg508_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1140_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg682_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg526_out;
SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg322_out;
SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg889_out;
SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg889_out;
SharedReg1163_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1163_out;
SharedReg1165_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1165_out;
SharedReg1137_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
SharedReg1142_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1142_out;
SharedReg525_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg525_out;
SharedReg76_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg76_out;
SharedReg1154_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1154_out;
SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg515_out;
SharedReg704_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg704_out;
SharedReg1139_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1139_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg505_out;
SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1135_out;
SharedReg699_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg699_out;
SharedReg726_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg726_out;
SharedReg1419_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1419_out;
SharedReg321_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg321_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg505_out;
SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg322_out;
SharedReg516_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg516_out;
SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1135_out;
SharedReg334_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg334_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg505_out;
SharedReg695_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg695_out;
SharedReg66_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg66_out;
SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1135_out;
SharedReg1149_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1149_out;
SharedReg893_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg893_out;
SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg330_out;
SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg330_out;
SharedReg712_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg712_out;
SharedReg1356_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1356_out;
SharedReg698_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg698_out;
SharedReg509_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg509_out;
SharedReg327_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg327_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg505_out;
SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg912_out;
SharedReg545_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg545_out;
SharedReg111_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg111_out;
SharedReg544_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg544_out;
SharedReg718_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg718_out;
SharedReg918_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg918_out;
SharedReg925_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg925_out;
SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg526_out;
SharedReg1347_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1347_out;
SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg526_out;
SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg526_out;
SharedReg533_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg533_out;
SharedReg713_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg713_out;
SharedReg99_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg99_out;
SharedReg950_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg950_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1142_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg525_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg76_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1154_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg515_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg704_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1139_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg699_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg726_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1419_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg321_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg516_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg334_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg695_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg66_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1135_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1149_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg889_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg893_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg330_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg712_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1356_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg698_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg509_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg327_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1163_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg545_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg111_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg544_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg718_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg918_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg925_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1347_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1165_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg533_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg713_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg99_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg950_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No52_out);

SharedReg715_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg715_out;
SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg883_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg1349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1349_out;
SharedReg529_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg529_out;
SharedReg1160_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1160_out;
SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1136_out;
SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
SharedReg702_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg702_out;
SharedReg706_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg706_out;
SharedReg78_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg78_out;
SharedReg1148_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1148_out;
SharedReg703_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg703_out;
SharedReg1144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1144_out;
SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg693_out;
SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg693_out;
SharedReg512_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg512_out;
SharedReg701_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg701_out;
SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1135_out;
SharedReg540_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg540_out;
SharedReg1350_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1350_out;
SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg93_out;
SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg694_out;
SharedReg339_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg339_out;
SharedReg522_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg522_out;
SharedReg698_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg698_out;
SharedReg319_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg319_out;
SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1139_out;
SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1135_out;
SharedReg323_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg323_out;
SharedReg1152_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1152_out;
SharedReg1137_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1137_out;
SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1347_out;
SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg317_out;
SharedReg67_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg67_out;
SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1139_out;
SharedReg891_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg891_out;
SharedReg1138_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1138_out;
SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1136_out;
Delay91No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast <= Delay91No1_out;
SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg694_out;
SharedReg1432_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1432_out;
SharedReg718_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg718_out;
SharedReg343_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg343_out;
SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg532_out;
SharedReg716_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg716_out;
SharedReg939_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg939_out;
SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1347_out;
SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1157_out;
SharedReg931_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg931_out;
SharedReg714_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg714_out;
SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1157_out;
SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg526_out;
SharedReg1162_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1162_out;
SharedReg120_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg120_out;
SharedReg1455_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1455_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg715_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg702_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg706_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg78_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1148_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg703_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1144_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg693_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg512_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg701_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg540_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1350_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg93_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg883_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg339_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg522_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg698_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg319_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1135_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg323_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1152_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1137_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1349_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg67_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1139_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg891_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1138_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => Delay91No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg694_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1432_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg529_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg718_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg343_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg716_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg939_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1347_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg931_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg714_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1157_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1160_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1162_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg120_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1455_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1136_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg554_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg733_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg733_out;
SharedReg347_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg347_out;
SharedReg1331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1331_out;
SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg547_out;
SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg348_out;
SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg100_out;
SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1354_out;
SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1354_out;
SharedReg1183_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1183_out;
SharedReg1185_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1185_out;
SharedReg1157_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1157_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg8_out;
SharedReg1162_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1162_out;
SharedReg546_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg546_out;
SharedReg105_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg105_out;
SharedReg1174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1174_out;
SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg10_out;
SharedReg724_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg724_out;
SharedReg1159_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1159_out;
SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg526_out;
SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg526_out;
SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1155_out;
SharedReg719_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg719_out;
SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg746_out;
SharedReg901_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg901_out;
SharedReg99_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg99_out;
SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg526_out;
SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg348_out;
SharedReg537_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg537_out;
SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1155_out;
SharedReg360_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg360_out;
SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg526_out;
SharedReg715_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg715_out;
SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg95_out;
SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1155_out;
SharedReg1169_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1169_out;
SharedReg921_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg921_out;
SharedReg356_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg356_out;
SharedReg373_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg373_out;
SharedReg555_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg555_out;
SharedReg940_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg940_out;
SharedReg951_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg951_out;
SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg380_out;
SharedReg124_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg124_out;
SharedReg950_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg950_out;
SharedReg381_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg381_out;
SharedReg752_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg752_out;
SharedReg1330_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1330_out;
SharedReg738_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg738_out;
SharedReg551_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg551_out;
SharedReg378_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg378_out;
SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg547_out;
SharedReg942_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg942_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1354_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1183_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1185_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1157_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1162_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg546_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg105_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg10_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg724_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1159_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg554_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg719_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg901_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg99_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg537_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg733_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg360_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg526_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg715_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg95_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1155_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1169_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg921_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg356_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg373_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg347_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg555_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg940_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg951_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg124_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg950_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg381_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg752_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1330_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg738_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg551_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg378_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg942_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg547_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg348_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No54_out);

SharedReg961_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg961_out;
SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg734_out;
SharedReg1177_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1177_out;
SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg547_out;
SharedReg1182_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1182_out;
SharedReg149_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg149_out;
SharedReg965_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg965_out;
SharedReg735_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg735_out;
SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg343_out;
SharedReg911_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg911_out;
SharedReg1430_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1430_out;
SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg550_out;
SharedReg1180_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1180_out;
SharedReg1156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1156_out;
SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg26_out;
SharedReg722_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg722_out;
SharedReg726_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg726_out;
SharedReg107_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg107_out;
SharedReg1168_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1168_out;
SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg28_out;
SharedReg1164_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1164_out;
SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg713_out;
SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg713_out;
SharedReg533_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg533_out;
SharedReg721_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg721_out;
SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1155_out;
SharedReg561_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg561_out;
SharedReg1431_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1431_out;
SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg338_out;
SharedReg714_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg714_out;
SharedReg122_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg122_out;
SharedReg543_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg543_out;
SharedReg718_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg718_out;
SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg345_out;
SharedReg1159_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1159_out;
SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1155_out;
SharedReg349_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg349_out;
SharedReg1172_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1172_out;
SharedReg1157_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1157_out;
SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1428_out;
SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg343_out;
SharedReg368_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg368_out;
SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg547_out;
SharedReg945_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg945_out;
SharedReg940_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg940_out;
SharedReg124_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg124_out;
SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg370_out;
SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1428_out;
SharedReg344_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg344_out;
SharedReg1179_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1179_out;
SharedReg949_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg949_out;
SharedReg1178_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1178_out;
SharedReg1176_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1176_out;
Delay91No3_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast <= Delay91No3_out;
SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg734_out;
SharedReg972_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg972_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg961_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg911_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1430_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1180_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1156_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1177_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg722_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg726_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1168_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg28_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1164_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg713_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg533_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg721_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg561_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1431_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg714_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg122_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg543_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1182_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg718_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1159_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1155_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg349_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1172_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1157_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg368_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg149_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg547_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg945_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg940_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg124_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1428_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg344_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1179_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg949_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1178_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg965_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1176_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => Delay91No3_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg734_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg972_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg735_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg343_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg772_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg772_out;
SharedReg977_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg977_out;
SharedReg758_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg758_out;
SharedReg572_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg572_out;
SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg164_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg568_out;
SharedReg1323_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1323_out;
SharedReg940_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg940_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg575_out;
SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg753_out;
SharedReg372_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg372_out;
SharedReg978_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg978_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg568_out;
SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg373_out;
SharedReg129_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg129_out;
SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1435_out;
SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1435_out;
SharedReg1203_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1203_out;
SharedReg1205_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1205_out;
SharedReg1177_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1177_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg11_out;
SharedReg570_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg570_out;
SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg8_out;
SharedReg1182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1182_out;
SharedReg567_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg567_out;
SharedReg134_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg134_out;
SharedReg1194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1194_out;
SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg10_out;
SharedReg744_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg744_out;
SharedReg1179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1179_out;
SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg547_out;
SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1175_out;
SharedReg739_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg739_out;
SharedReg766_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg766_out;
SharedReg929_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg929_out;
SharedReg128_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg128_out;
SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg547_out;
SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg373_out;
SharedReg558_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg558_out;
SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1175_out;
SharedReg386_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg386_out;
SharedReg1338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1338_out;
SharedReg1001_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1001_out;
SharedReg970_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg970_out;
SharedReg143_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg143_out;
SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg753_out;
SharedReg1208_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1208_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg568_out;
SharedReg755_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg755_out;
SharedReg368_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg368_out;
SharedReg1195_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1195_out;
SharedReg1209_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1209_out;
SharedReg979_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg979_out;
SharedReg409_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg409_out;
SharedReg188_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg188_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg772_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg977_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg372_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg978_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg129_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1435_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1203_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg758_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1205_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1177_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg570_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg572_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg567_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg134_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg10_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg744_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg164_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg739_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg766_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg929_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg128_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg547_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg373_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg558_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1175_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg386_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1001_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg970_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg143_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg753_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1208_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg755_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg368_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1195_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1323_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1209_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg979_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg409_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg188_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg940_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No56_out);

SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1199_out;
SharedReg1330_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1330_out;
SharedReg1198_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1198_out;
SharedReg1196_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1196_out;
Delay91No4_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= Delay91No4_out;
SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg754_out;
SharedReg1002_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1002_out;
SharedReg991_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg991_out;
SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg754_out;
SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1197_out;
SharedReg568_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg568_out;
SharedReg1202_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1202_out;
SharedReg391_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg391_out;
SharedReg995_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg995_out;
SharedReg755_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg755_out;
SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg368_out;
SharedReg941_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg941_out;
SharedReg1323_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1323_out;
SharedReg571_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg571_out;
SharedReg1200_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1200_out;
SharedReg1176_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1176_out;
SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg29_out;
SharedReg753_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg753_out;
SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg26_out;
SharedReg742_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg742_out;
SharedReg746_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg746_out;
SharedReg136_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg136_out;
SharedReg1188_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1188_out;
SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg28_out;
SharedReg1184_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1184_out;
SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg733_out;
SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg733_out;
SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg554_out;
SharedReg741_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg741_out;
SharedReg1175_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1175_out;
SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg582_out;
SharedReg1324_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1324_out;
SharedReg121_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg121_out;
SharedReg734_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg734_out;
SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg364_out;
SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg564_out;
SharedReg738_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg738_out;
SharedReg370_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg370_out;
SharedReg971_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg971_out;
SharedReg963_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg963_out;
SharedReg1344_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1344_out;
SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg161_out;
SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1195_out;
SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg581_out;
SharedReg760_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg760_out;
SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1199_out;
SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1195_out;
SharedReg402_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg402_out;
SharedReg1212_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1212_out;
SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1197_out;
SharedReg1321_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1321_out;
SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg368_out;
SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg396_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1330_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg568_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1202_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg391_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg995_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg755_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg941_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1323_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg571_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1198_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1200_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1176_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg753_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1196_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg742_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg746_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg136_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1188_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg28_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1184_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg733_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg741_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => Delay91No4_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1175_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1324_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg121_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg734_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg364_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg738_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg370_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg971_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg963_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1344_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg760_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1199_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1195_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg402_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1212_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1002_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1321_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg368_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg991_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg754_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1197_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg775_out;
SharedReg154_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1215_out;
SharedReg1229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1229_out;
SharedReg1009_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1009_out;
SharedReg195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg195_out;
SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg431_out;
SharedReg792_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg792_out;
SharedReg1007_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1007_out;
SharedReg778_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg778_out;
SharedReg593_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg593_out;
SharedReg406_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg589_out;
SharedReg1000_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1000_out;
SharedReg968_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg968_out;
SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg589_out;
SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg589_out;
SharedReg596_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg596_out;
SharedReg773_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg773_out;
SharedReg400_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg400_out;
SharedReg1036_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1036_out;
SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg589_out;
SharedReg401_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg401_out;
SharedReg159_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg159_out;
SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1328_out;
SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1328_out;
SharedReg1223_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1223_out;
SharedReg793_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg793_out;
SharedReg1197_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1197_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg11_out;
SharedReg591_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg591_out;
SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg8_out;
SharedReg1202_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1202_out;
SharedReg588_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg588_out;
SharedReg165_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg165_out;
SharedReg1214_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1214_out;
SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg10_out;
SharedReg764_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg764_out;
SharedReg1199_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1199_out;
SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg568_out;
SharedReg1195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1195_out;
SharedReg759_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg759_out;
SharedReg786_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg786_out;
SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg775_out;
SharedReg426_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg426_out;
SharedReg1028_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1028_out;
SharedReg1027_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1027_out;
SharedReg1374_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1374_out;
SharedReg595_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg595_out;
SharedReg429_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg429_out;
SharedReg987_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg987_out;
SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg187_out;
SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg589_out;
SharedReg188_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg188_out;
SharedReg600_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg600_out;
SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1215_out;
SharedReg444_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg444_out;
SharedReg1392_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1392_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg593_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1000_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg968_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg596_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg773_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg400_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1036_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg401_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg159_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1328_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1223_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg793_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1197_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg591_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1202_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg588_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg165_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1009_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1214_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg10_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg764_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1199_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg759_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg786_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg775_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg195_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg426_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1028_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1027_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1374_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg595_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg429_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg987_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg589_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg188_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg600_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1215_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg444_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1392_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg792_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1007_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg778_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No58_out);

SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1215_out;
SharedReg189_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg1232_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1232_out;
SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1217_out;
SharedReg968_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg968_out;
SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg426_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg1219_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1219_out;
SharedReg977_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg977_out;
SharedReg1218_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1218_out;
SharedReg1216_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1216_out;
Delay91No5_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= Delay91No5_out;
SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg774_out;
SharedReg1377_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1377_out;
SharedReg1050_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1050_out;
SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg774_out;
SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1217_out;
SharedReg589_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg589_out;
SharedReg1222_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1222_out;
SharedReg421_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg421_out;
SharedReg1054_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1054_out;
SharedReg775_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg775_out;
SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg396_out;
SharedReg969_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg969_out;
SharedReg1000_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1000_out;
SharedReg592_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg592_out;
SharedReg1235_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1235_out;
SharedReg1196_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1196_out;
SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg29_out;
SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg773_out;
SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg26_out;
SharedReg762_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg762_out;
SharedReg766_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg766_out;
SharedReg167_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg167_out;
SharedReg1208_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1208_out;
SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg28_out;
SharedReg1204_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1204_out;
SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg753_out;
SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg753_out;
SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg575_out;
SharedReg761_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg761_out;
SharedReg1195_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1195_out;
SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg603_out;
SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1215_out;
SharedReg198_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg198_out;
SharedReg1041_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1041_out;
SharedReg1055_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1055_out;
SharedReg1398_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1398_out;
SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg773_out;
SharedReg455_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg455_out;
SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1030_out;
SharedReg181_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg181_out;
SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg774_out;
SharedReg422_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg422_out;
SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg606_out;
SharedReg778_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg778_out;
SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg185_out;
SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1030_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1216_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay91No5_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1377_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1050_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg589_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1222_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg421_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1232_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1054_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg775_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg969_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1000_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg592_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1235_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1196_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1217_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg762_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg766_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg167_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg968_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1208_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg28_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1204_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg753_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg761_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1195_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1215_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg198_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1041_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1055_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1398_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg773_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg455_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg181_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg774_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg422_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg426_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg778_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1030_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1219_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg977_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1218_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add11_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_5_impl_out,
                 X => Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast);

SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg430_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg610_out;
SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg431_out;
SharedReg621_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg621_out;
SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1235_out;
SharedReg253_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg253_out;
SharedReg1312_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1312_out;
SharedReg795_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg183_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg183_out;
SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1235_out;
SharedReg1249_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1249_out;
SharedReg1037_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1037_out;
SharedReg439_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg439_out;
SharedReg240_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg240_out;
SharedReg812_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg812_out;
SharedReg1382_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1382_out;
SharedReg798_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg798_out;
SharedReg614_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg614_out;
SharedReg436_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg436_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg610_out;
SharedReg1375_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1375_out;
SharedReg1027_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1027_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg610_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg610_out;
SharedReg617_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg617_out;
SharedReg793_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg793_out;
SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg430_out;
SharedReg631_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg631_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg610_out;
SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg431_out;
SharedReg188_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg188_out;
SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1005_out;
SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1005_out;
SharedReg1243_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1243_out;
SharedReg813_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg813_out;
SharedReg1217_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1217_out;
SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg11_out;
SharedReg612_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg612_out;
SharedReg16_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg8_out;
SharedReg1222_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1222_out;
SharedReg609_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg609_out;
SharedReg193_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg193_out;
SharedReg1234_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1234_out;
SharedReg10_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg13_out;
SharedReg613_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg613_out;
SharedReg1044_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1044_out;
SharedReg1067_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1067_out;
SharedReg811_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg811_out;
SharedReg620_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg620_out;
SharedReg804_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg804_out;
SharedReg1239_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1239_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg610_out;
SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg610_out;
SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1235_out;
SharedReg799_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg799_out;
SharedReg826_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg826_out;
SharedReg815_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg815_out;
   MUX_Add11_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1249_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1037_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg439_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg240_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg812_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1382_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg798_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg614_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg436_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1375_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1027_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg617_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg793_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg430_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg631_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg431_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg621_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg188_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1005_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1243_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg813_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1217_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg3_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg17_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg11_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg612_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg16_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg8_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1222_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg609_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg193_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1234_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg10_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg253_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg13_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg613_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1044_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1067_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg811_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg620_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg804_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1239_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg610_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1312_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg799_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg826_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg815_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg795_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg183_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1235_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_5_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_0_out,
                 Y => Delay1No60_out);

SharedReg208_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg794_out;
SharedReg451_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg627_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg627_out;
SharedReg798_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg798_out;
SharedReg428_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg428_out;
SharedReg1376_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1376_out;
SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1235_out;
SharedReg432_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg432_out;
SharedReg1252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1252_out;
SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1237_out;
SharedReg1027_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1027_out;
SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg426_out;
SharedReg235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg235_out;
SharedReg1239_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1239_out;
SharedReg1035_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1035_out;
SharedReg1238_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1238_out;
SharedReg1236_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1236_out;
Delay91No6_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast <= Delay91No6_out;
SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg794_out;
SharedReg1299_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1299_out;
SharedReg1079_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1079_out;
SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg794_out;
SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1237_out;
SharedReg610_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg610_out;
SharedReg1242_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1242_out;
SharedReg450_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg450_out;
SharedReg1257_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1257_out;
SharedReg795_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg795_out;
SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg426_out;
SharedReg1028_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1028_out;
SharedReg1375_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1375_out;
SharedReg613_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg613_out;
SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1255_out;
SharedReg1216_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1216_out;
SharedReg19_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg29_out;
SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg793_out;
SharedReg34_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg26_out;
SharedReg782_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg782_out;
SharedReg786_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg786_out;
SharedReg195_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg195_out;
SharedReg1228_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1228_out;
SharedReg28_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg31_out;
SharedReg797_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg797_out;
SharedReg1386_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1386_out;
SharedReg1069_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1069_out;
SharedReg622_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg622_out;
SharedReg803_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg803_out;
SharedReg1244_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1244_out;
SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg793_out;
SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg793_out;
SharedReg617_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg617_out;
SharedReg801_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg801_out;
SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1235_out;
SharedReg645_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg645_out;
SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1255_out;
   MUX_Add11_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1027_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1239_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1035_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1238_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1236_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay91No6_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg451_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1299_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1079_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg794_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1237_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg610_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1242_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg450_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1257_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg795_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg627_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg426_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1028_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1375_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg613_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1216_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg19_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg35_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg33_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg798_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg29_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg34_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg26_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg782_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg786_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg195_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1228_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg28_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg27_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg428_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg797_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1386_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1069_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg622_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg803_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1244_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg793_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg617_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1376_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg801_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg645_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1255_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1235_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg432_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_5_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add11_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_8_impl_out,
                 X => Delay1No62_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg15_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg16_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg17_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg469_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg469_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg652_out;
SharedReg1097_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1097_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg652_out;
SharedReg261_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg261_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg652_out;
SharedReg240_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg240_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg652_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg652_out;
SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg467_out;
SharedReg668_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg668_out;
SharedReg1302_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1302_out;
SharedReg654_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg654_out;
SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg461_out;
SharedReg659_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg659_out;
SharedReg672_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg672_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg652_out;
SharedReg1093_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1093_out;
SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg833_out;
SharedReg1474_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1474_out;
SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg467_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg652_out;
SharedReg1096_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1096_out;
SharedReg1278_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1278_out;
SharedReg1285_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1285_out;
SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg652_out;
SharedReg265_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg265_out;
SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg833_out;
SharedReg466_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg466_out;
SharedReg663_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg663_out;
SharedReg852_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg852_out;
SharedReg838_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg838_out;
SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1275_out;
SharedReg1086_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1086_out;
SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg461_out;
SharedReg844_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg844_out;
SharedReg656_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg656_out;
SharedReg1282_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1282_out;
SharedReg1277_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1277_out;
SharedReg835_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg835_out;
SharedReg1289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1289_out;
SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1275_out;
SharedReg1279_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1279_out;
SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1275_out;
SharedReg1464_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1464_out;
   MUX_Add11_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg261_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg240_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg668_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1302_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg654_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg8_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg659_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg672_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1093_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1474_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg467_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1096_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1278_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg15_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1285_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg265_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg833_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg466_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg663_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg852_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg838_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1086_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg16_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg461_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg844_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg656_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1282_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1277_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg835_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1279_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1275_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg17_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1464_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg469_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1097_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg652_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add11_8_impl_0_LUT_out,
                 oMux => MUX_Add11_8_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_8_impl_0_out,
                 Y => Delay1No62_out);

SharedReg19_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg33_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg33_out;
SharedReg34_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg35_out;
SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg834_out;
SharedReg659_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg659_out;
SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg833_out;
SharedReg1095_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1095_out;
SharedReg267_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg267_out;
SharedReg835_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg835_out;
SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg834_out;
SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg838_out;
SharedReg469_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg469_out;
SharedReg837_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg837_out;
SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg457_out;
SharedReg652_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg652_out;
SharedReg1087_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1087_out;
SharedReg846_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg846_out;
SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1277_out;
SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1275_out;
SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1277_out;
SharedReg1089_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1089_out;
SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1280_out;
SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg457_out;
SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1280_out;
SharedReg1086_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1086_out;
SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1279_out;
SharedReg1459_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1459_out;
SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg457_out;
SharedReg1282_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1282_out;
SharedReg286_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg286_out;
SharedReg669_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg669_out;
Delay91No8_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_35_cast <= Delay91No8_out;
SharedReg1278_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1278_out;
SharedReg480_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg480_out;
SharedReg1292_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1292_out;
SharedReg1108_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1108_out;
SharedReg262_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg262_out;
SharedReg1457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1457_out;
SharedReg1284_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1284_out;
SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1279_out;
SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1276_out;
SharedReg842_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg842_out;
SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1276_out;
SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1275_out;
SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg838_out;
SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1277_out;
SharedReg841_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg841_out;
SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg833_out;
   MUX_Add11_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg267_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg835_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg469_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg837_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg652_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1087_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg846_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg26_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1089_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1280_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1086_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1459_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg33_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1282_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg286_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg669_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay91No8_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1278_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg480_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1292_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1108_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg262_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg34_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1457_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1284_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1279_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg842_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1276_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1275_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg838_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1277_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg841_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg35_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg834_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg659_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg833_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1095_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add11_8_impl_1_LUT_out,
                 oMux => MUX_Add11_8_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_8_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No64_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1535_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1482_out;
SharedReg1400_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1400_out;
SharedReg1588_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1634_out;
SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg856_out;
SharedReg1486_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1487_out;
SharedReg1405_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1405_out;
SharedReg1489_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1604_out;
SharedReg860_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg860_out;
SharedReg1600_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1600_out;
SharedReg1411_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1411_out;
SharedReg1631_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1548_out;
SharedReg1412_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1412_out;
SharedReg1524_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1635_out;
SharedReg45_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg45_out;
SharedReg1527_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1621_out;
SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg48_out;
SharedReg1517_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1534_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1535_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1521_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1634_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg856_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1486_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1487_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1405_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1489_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1630_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1490_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1603_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1604_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1522_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg860_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1600_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1411_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1631_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1495_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1548_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1412_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1524_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1641_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1635_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1585_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg45_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1527_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1528_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1498_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1499_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1500_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1501_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1502_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1591_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1503_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1536_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1504_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1593_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1556_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1506_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1507_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1508_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1509_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1510_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1560_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1511_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1523_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1512_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1513_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1565_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1621_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1517_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1518_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1519_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1520_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1537_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1610_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1532_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1582_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1534_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1482_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1400_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1588_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No64_out);

SharedReg1422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1422_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg1424_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1424_out;
SharedReg60_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg36_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg37_out;
SharedReg1648_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1648_out;
SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1400_out;
SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg1640_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1640_out;
SharedReg295_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg295_out;
SharedReg297_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg297_out;
SharedReg1594_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1594_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg44_out;
SharedReg1406_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1406_out;
SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg42_out;
SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg859_out;
SharedReg861_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg861_out;
SharedReg1601_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1601_out;
SharedReg864_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg864_out;
SharedReg1633_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1633_out;
SharedReg1412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1412_out;
SharedReg301_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg301_out;
SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg48_out;
SharedReg1628_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1628_out;
SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg47_out;
SharedReg1415_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1415_out;
SharedReg1416_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1416_out;
SharedReg1576_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1576_out;
SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg46_out;
SharedReg866_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg866_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg36_out;
SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1400_out;
SharedReg290_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg290_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg36_out;
SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1401_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg36_out;
SharedReg291_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg291_out;
SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1401_out;
SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg43_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg44_out;
SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg296_out;
SharedReg1407_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1407_out;
SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg296_out;
SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg43_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg44_out;
SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg39_out;
SharedReg298_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg298_out;
SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg39_out;
SharedReg1410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1410_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg37_out;
SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg859_out;
SharedReg1566_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1566_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg36_out;
SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg855_out;
SharedReg58_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg58_out;
SharedReg311_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg311_out;
SharedReg59_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg59_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1640_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg295_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg297_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1594_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1406_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg861_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1601_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg864_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1633_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1412_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg301_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1628_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg47_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1415_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1416_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1424_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1576_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg866_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg290_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg60_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg291_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1401_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1407_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg296_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg298_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1410_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg859_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1566_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg855_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg58_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg311_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg59_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1648_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1400_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No66_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1518_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1482_out;
SharedReg1347_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1347_out;
SharedReg1588_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1634_out;
SharedReg885_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg885_out;
SharedReg1486_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1487_out;
SharedReg1352_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1352_out;
SharedReg1489_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1604_out;
SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg889_out;
SharedReg1600_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1600_out;
SharedReg1358_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1358_out;
SharedReg1631_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1548_out;
SharedReg1359_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1359_out;
SharedReg1524_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1635_out;
SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg75_out;
SharedReg1527_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1621_out;
SharedReg78_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg78_out;
SharedReg1517_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1517_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1518_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1519_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1585_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1536_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1523_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1537_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1482_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1347_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1588_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1634_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg885_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1486_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1520_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1487_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1352_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1489_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1630_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1490_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1603_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1604_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg889_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1600_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1358_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1610_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1631_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1495_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1548_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1359_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1524_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1641_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1635_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1527_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1532_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1498_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1500_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1501_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1502_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1591_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1503_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1504_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1593_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1556_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1582_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1506_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1507_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1508_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1509_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1510_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1560_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1511_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1512_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1513_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1514_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1534_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1565_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1621_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg78_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1517_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1535_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1521_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1522_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No66_out);

SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg1402_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1402_out;
SharedReg311_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg311_out;
SharedReg336_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg336_out;
SharedReg88_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg1367_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1367_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg66_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg66_out;
SharedReg1369_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1369_out;
SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg66_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg66_out;
SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg67_out;
SharedReg1648_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1648_out;
SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1347_out;
SharedReg884_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg884_out;
SharedReg1640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1640_out;
SharedReg322_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg322_out;
SharedReg324_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg324_out;
SharedReg1594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1594_out;
SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg74_out;
SharedReg1353_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1353_out;
SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg72_out;
SharedReg888_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg888_out;
SharedReg890_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg890_out;
SharedReg1601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1601_out;
SharedReg893_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg893_out;
SharedReg1633_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1633_out;
SharedReg1359_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1359_out;
SharedReg328_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg328_out;
SharedReg78_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg78_out;
SharedReg1628_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1628_out;
SharedReg77_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg77_out;
SharedReg1362_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1362_out;
SharedReg1363_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1363_out;
SharedReg1576_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1576_out;
SharedReg76_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg76_out;
SharedReg895_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg895_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg66_out;
SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1347_out;
SharedReg317_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg317_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg66_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg66_out;
SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1348_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg66_out;
SharedReg318_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg318_out;
SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1348_out;
SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg73_out;
SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg74_out;
SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg323_out;
SharedReg1354_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1354_out;
SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg323_out;
SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg73_out;
SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg74_out;
SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg69_out;
SharedReg325_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg325_out;
SharedReg293_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg293_out;
SharedReg1357_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1357_out;
SharedReg291_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg291_out;
SharedReg1406_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1406_out;
SharedReg1566_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1566_out;
SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg290_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1369_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1648_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg884_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg322_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg324_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1353_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg888_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg890_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg893_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1633_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1402_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1359_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg328_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg78_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1628_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg77_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1362_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1363_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1576_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg76_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg895_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg311_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1347_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg317_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg318_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1348_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg336_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1354_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg323_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg73_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg325_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg293_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1357_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg291_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1406_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1566_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg290_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1367_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No68_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1512_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1621_out;
SharedReg330_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg330_out;
SharedReg1517_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1482_out;
SharedReg1428_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1428_out;
SharedReg1588_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1634_out;
SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg913_out;
SharedReg1486_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1487_out;
SharedReg1433_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1433_out;
SharedReg1489_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1604_out;
SharedReg917_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg917_out;
SharedReg1600_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1600_out;
SharedReg1439_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1439_out;
SharedReg1631_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1548_out;
SharedReg1440_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1440_out;
SharedReg1524_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1635_out;
SharedReg104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg104_out;
SharedReg1527_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1511_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1512_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1513_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1610_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1532_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1582_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1534_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1535_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1521_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1522_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1585_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1536_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1523_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1514_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1537_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1482_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1428_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1588_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1634_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1486_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1487_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1433_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1489_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1565_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1630_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1490_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1603_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1604_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg917_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1600_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1439_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1631_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1548_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1621_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1440_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1524_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1641_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1635_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1527_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1528_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1498_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1499_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1500_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg330_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1501_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1502_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1591_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1503_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1504_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1593_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1556_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1507_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1508_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1517_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1509_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1510_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1560_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1511_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1518_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1519_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1520_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No68_out);

SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg69_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg920_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg67_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg67_out;
SharedReg888_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg888_out;
SharedReg1566_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1566_out;
SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg1349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1349_out;
SharedReg336_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg336_out;
SharedReg362_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg362_out;
SharedReg116_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg116_out;
SharedReg1448_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1448_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg1450_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1450_out;
SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg117_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg95_out;
SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg96_out;
SharedReg1648_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1648_out;
SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1428_out;
SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg912_out;
SharedReg1640_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1640_out;
SharedReg348_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg348_out;
SharedReg350_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg350_out;
SharedReg1594_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1594_out;
SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg103_out;
SharedReg1434_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1434_out;
SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg101_out;
SharedReg916_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg916_out;
SharedReg918_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg918_out;
SharedReg1601_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1601_out;
SharedReg921_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg921_out;
SharedReg1633_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1633_out;
SharedReg1440_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1440_out;
SharedReg354_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg354_out;
SharedReg107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg107_out;
SharedReg1628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1628_out;
SharedReg106_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg106_out;
SharedReg1443_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1443_out;
SharedReg1444_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1444_out;
SharedReg1576_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1576_out;
SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg105_out;
SharedReg923_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg923_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg95_out;
SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1428_out;
SharedReg343_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg343_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg95_out;
SharedReg1429_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1429_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg95_out;
SharedReg344_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg344_out;
SharedReg911_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg911_out;
SharedReg102_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg102_out;
SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg103_out;
SharedReg349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg349_out;
SharedReg1435_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1435_out;
SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg101_out;
SharedReg324_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg324_out;
SharedReg325_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg325_out;
SharedReg320_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg320_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg336_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg362_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg116_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1448_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1450_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1648_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1640_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg348_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg350_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1594_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg67_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1434_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg916_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg918_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1601_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg921_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1633_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1440_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg354_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg888_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg106_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1443_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1444_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1576_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg923_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1428_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg343_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1566_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1429_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg344_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg911_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg102_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg349_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1435_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg324_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg325_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg320_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No70_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1506_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1621_out;
SharedReg107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg107_out;
SharedReg1517_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1482_out;
SharedReg1321_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1321_out;
SharedReg1588_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1634_out;
SharedReg943_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg943_out;
SharedReg1486_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1487_out;
SharedReg1326_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1326_out;
SharedReg1489_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1604_out;
SharedReg947_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg947_out;
SharedReg1600_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1600_out;
SharedReg1332_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1332_out;
SharedReg1631_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1548_out;
SharedReg1333_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1333_out;
SharedReg1524_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1635_out;
SharedReg133_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg133_out;
SharedReg1527_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1556_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1506_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1507_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1565_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1621_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1517_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1518_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1519_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1520_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1610_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1532_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1582_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1508_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1534_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1535_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1521_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1522_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1585_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1536_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1523_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1537_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1482_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1321_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1509_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1588_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1634_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg943_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1486_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1487_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1326_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1489_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1630_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1490_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1603_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1510_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1604_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg947_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1600_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1332_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1631_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1495_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1548_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1333_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1524_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1641_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1560_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1635_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg133_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1527_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1528_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1498_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1499_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1500_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1501_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1502_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1591_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1511_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1503_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1504_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1593_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1512_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1514_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No70_out);

SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg947_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg947_out;
SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg349_out;
SharedReg102_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg102_out;
SharedReg103_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg103_out;
SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg98_out;
SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg351_out;
SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg98_out;
SharedReg1438_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1438_out;
SharedReg96_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg916_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg916_out;
SharedReg1566_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1566_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg343_out;
SharedReg1430_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1430_out;
SharedReg362_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg362_out;
SharedReg388_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg388_out;
SharedReg145_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg145_out;
SharedReg1341_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1341_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg124_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg124_out;
SharedReg1343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1343_out;
SharedReg146_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg146_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg124_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg124_out;
SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg125_out;
SharedReg1648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1648_out;
SharedReg1321_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1321_out;
SharedReg942_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg942_out;
SharedReg1640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1640_out;
SharedReg373_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg373_out;
SharedReg375_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg375_out;
SharedReg1594_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1594_out;
SharedReg132_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg132_out;
SharedReg1327_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1327_out;
SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg349_out;
SharedReg946_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg946_out;
SharedReg948_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg948_out;
SharedReg1601_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1601_out;
SharedReg951_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg951_out;
SharedReg1633_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1633_out;
SharedReg1333_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1333_out;
SharedReg379_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg379_out;
SharedReg136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg136_out;
SharedReg1628_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1628_out;
SharedReg135_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg135_out;
SharedReg1336_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1336_out;
SharedReg1337_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1337_out;
SharedReg1576_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1576_out;
SharedReg134_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg134_out;
SharedReg953_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg953_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg343_out;
SharedReg940_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg940_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg124_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg343_out;
SharedReg941_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg941_out;
SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg343_out;
SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg125_out;
SharedReg1429_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1429_out;
SharedReg350_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg350_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg916_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1566_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1430_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg362_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg388_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg947_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg145_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1341_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg146_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1321_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg942_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg373_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg375_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1594_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg132_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1327_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg349_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg946_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg102_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg948_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1601_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg951_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1633_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1333_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg379_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1628_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg135_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1336_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg103_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1337_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1576_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg134_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg953_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg940_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg941_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg343_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1429_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg350_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg351_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg98_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1438_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No72_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1501_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1621_out;
SharedReg136_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg136_out;
SharedReg1517_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1482_out;
SharedReg998_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg998_out;
SharedReg1588_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1634_out;
SharedReg971_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg971_out;
SharedReg1486_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1487_out;
SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1003_out;
SharedReg1489_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1604_out;
SharedReg975_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg975_out;
SharedReg1600_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1600_out;
SharedReg1009_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1009_out;
SharedReg1631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1548_out;
SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1010_out;
SharedReg1524_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1635_out;
SharedReg164_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg164_out;
SharedReg1527_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1500_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1501_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1502_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1509_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1510_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1560_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1511_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1512_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1513_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1514_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1565_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1621_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg136_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1591_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1517_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1519_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1520_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1610_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1532_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1582_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1534_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1535_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1521_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1503_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1522_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1585_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1536_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1523_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1537_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1482_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg998_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1588_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1634_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg971_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1504_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1486_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1487_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1489_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1490_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1603_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1604_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg975_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1600_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1593_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1009_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1495_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1548_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1524_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1641_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1635_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg164_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1527_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1556_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1528_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1498_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1499_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1500_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1506_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1507_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1508_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No72_out);

SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg124_out;
SharedReg1322_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1322_out;
SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg369_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg369_out;
SharedReg941_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg941_out;
SharedReg131_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg131_out;
SharedReg132_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg132_out;
SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg374_out;
SharedReg1328_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1328_out;
SharedReg130_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg130_out;
SharedReg350_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg350_out;
SharedReg351_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg351_out;
SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
SharedReg376_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg376_out;
SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg127_out;
SharedReg1331_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1331_out;
SharedReg125_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg125_out;
SharedReg946_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg946_out;
SharedReg1566_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1566_out;
SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg368_out;
SharedReg1323_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1323_out;
SharedReg388_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg388_out;
SharedReg176_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg176_out;
SharedReg389_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg389_out;
SharedReg989_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg989_out;
SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg154_out;
SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg154_out;
SharedReg992_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg992_out;
SharedReg390_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg390_out;
SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg154_out;
SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg154_out;
SharedReg155_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg155_out;
SharedReg1648_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1648_out;
SharedReg998_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg998_out;
SharedReg970_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg970_out;
SharedReg1640_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1640_out;
SharedReg401_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg401_out;
SharedReg403_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg403_out;
SharedReg1594_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1594_out;
SharedReg162_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg162_out;
SharedReg1004_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1004_out;
SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg374_out;
SharedReg974_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg974_out;
SharedReg976_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg976_out;
SharedReg1601_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1601_out;
SharedReg979_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg979_out;
SharedReg1633_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1633_out;
SharedReg1010_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1010_out;
SharedReg407_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg407_out;
SharedReg167_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg167_out;
SharedReg1628_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1628_out;
SharedReg166_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg166_out;
SharedReg1013_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1013_out;
SharedReg1014_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1014_out;
SharedReg1576_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1576_out;
SharedReg165_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg165_out;
SharedReg981_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg981_out;
SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg124_out;
SharedReg1321_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1321_out;
SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg368_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg130_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg350_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg351_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg376_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg127_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1331_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg125_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg946_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1566_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1322_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1323_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg388_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg176_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg389_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg989_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg992_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg390_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg154_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg155_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1648_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg998_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg970_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1640_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg369_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg401_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg403_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1594_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg162_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1004_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg974_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg976_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1601_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg979_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg941_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1633_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1010_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg407_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg167_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1628_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg166_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1013_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1014_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1576_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg165_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg131_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg981_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg124_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1321_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg368_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg132_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg374_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1328_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product4_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_5_impl_out,
                 X => Delay1No74_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1635_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1635_out;
SharedReg406_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg406_out;
SharedReg1527_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1621_out;
SharedReg167_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg167_out;
SharedReg1517_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1482_out;
SharedReg1373_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1373_out;
SharedReg1588_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1634_out;
SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1030_out;
SharedReg1486_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1487_out;
SharedReg1378_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1378_out;
SharedReg1489_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1604_out;
SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1033_out;
SharedReg1600_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1600_out;
SharedReg1384_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1384_out;
SharedReg1631_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1548_out;
SharedReg1385_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1385_out;
SharedReg1524_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1641_out;
   MUX_Product4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1635_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg406_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1503_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1504_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1593_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1556_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1506_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1507_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1508_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1509_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1510_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1560_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1527_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1511_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1512_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1513_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1514_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1565_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1621_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg167_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1517_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1518_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1519_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1528_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1520_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1610_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1532_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1582_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1534_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1535_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1521_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1522_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1585_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1536_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1498_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1523_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1537_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1482_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1373_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1588_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1634_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1486_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1487_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1378_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1499_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1489_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1630_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1490_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1603_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1604_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1600_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1384_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1631_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1495_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1500_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1548_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1385_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1524_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1641_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1501_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1502_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1591_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_5_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_0_out,
                 Y => Delay1No74_out);

SharedReg1389_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1389_out;
SharedReg1576_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1576_out;
SharedReg407_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg407_out;
SharedReg1040_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1040_out;
SharedReg368_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg998_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg396_out;
SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg154_out;
SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg154_out;
SharedReg999_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg999_out;
SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg154_out;
SharedReg397_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg397_out;
SharedReg969_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg969_out;
SharedReg161_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg161_out;
SharedReg162_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg162_out;
SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg402_out;
SharedReg1005_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1005_out;
SharedReg160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg160_out;
SharedReg375_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg375_out;
SharedReg376_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg376_out;
SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg157_out;
SharedReg404_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg404_out;
SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg157_out;
SharedReg1008_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1008_out;
SharedReg155_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg155_out;
SharedReg974_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg974_out;
SharedReg1566_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1566_out;
SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg396_out;
SharedReg1000_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1000_out;
SharedReg176_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg176_out;
SharedReg419_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg419_out;
SharedReg177_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg177_out;
SharedReg1021_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1021_out;
SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg183_out;
SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg183_out;
SharedReg1023_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1023_out;
SharedReg178_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg178_out;
SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg183_out;
SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg183_out;
SharedReg184_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg184_out;
SharedReg1648_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1648_out;
SharedReg1373_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1373_out;
SharedReg1029_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1029_out;
SharedReg1640_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1640_out;
SharedReg431_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg431_out;
SharedReg433_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg433_out;
SharedReg1594_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1594_out;
SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg191_out;
SharedReg1379_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1379_out;
SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg402_out;
SharedReg1032_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1032_out;
SharedReg1034_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1034_out;
SharedReg1601_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1601_out;
SharedReg1037_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1037_out;
SharedReg1633_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1633_out;
SharedReg1385_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1385_out;
SharedReg437_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg437_out;
SharedReg195_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg195_out;
SharedReg1628_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1628_out;
SharedReg194_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg194_out;
SharedReg1388_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1388_out;
   MUX_Product4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1389_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1576_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg397_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg969_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg161_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg162_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1005_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg375_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg376_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg407_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg404_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg157_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1008_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg155_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg974_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1566_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1040_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1000_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg176_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg419_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg177_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1021_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1023_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg178_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg368_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg183_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg184_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1648_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1373_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1029_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1640_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg431_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg433_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1594_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg998_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1379_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg402_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1032_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1034_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1601_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1037_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1633_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1385_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg437_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg396_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg195_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1628_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg194_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1388_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg154_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg999_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_5_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product4_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_6_impl_out,
                 X => Delay1No76_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1067_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1067_out;
SharedReg1631_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1548_out;
SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1068_out;
SharedReg1524_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1635_out;
SharedReg192_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg192_out;
SharedReg1527_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1621_out;
SharedReg195_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg195_out;
SharedReg1517_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1482_out;
SharedReg1295_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1295_out;
SharedReg1588_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1634_out;
SharedReg1060_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1060_out;
SharedReg1486_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1487_out;
SharedReg1300_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1300_out;
SharedReg1489_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1604_out;
SharedReg1380_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1380_out;
SharedReg1600_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1600_out;
   MUX_Product4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1067_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1631_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1528_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1498_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1499_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1500_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1501_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1502_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1591_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1503_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1504_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1593_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1495_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1556_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1506_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1507_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1508_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1509_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1510_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1560_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1511_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1512_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1513_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1548_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1514_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1565_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1621_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg195_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1517_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1518_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1519_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1520_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1610_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1532_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1582_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1534_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1535_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1521_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1522_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1585_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1536_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1523_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1537_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1482_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1524_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1295_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1588_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1634_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1060_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1486_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1487_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1300_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1489_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1630_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1490_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1641_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1603_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1604_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1380_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1600_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1635_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg192_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1527_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_6_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_0_out,
                 Y => Delay1No76_out);

SharedReg1633_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1633_out;
SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1068_out;
SharedReg220_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg439_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg1628_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1628_out;
SharedReg438_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
SharedReg1071_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1071_out;
SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1072_out;
SharedReg1576_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1576_out;
SharedReg193_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg193_out;
SharedReg1389_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1389_out;
SharedReg396_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg396_out;
SharedReg1373_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1373_out;
SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg426_out;
SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg183_out;
SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg183_out;
SharedReg1374_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1374_out;
SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg183_out;
SharedReg427_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg427_out;
SharedReg1028_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1028_out;
SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg190_out;
SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg191_out;
SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg432_out;
SharedReg1380_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1380_out;
SharedReg189_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg189_out;
SharedReg403_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg403_out;
SharedReg404_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg404_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg186_out;
SharedReg434_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg434_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg186_out;
SharedReg1383_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1383_out;
SharedReg184_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg184_out;
SharedReg1032_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1032_out;
SharedReg1566_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1566_out;
SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg426_out;
SharedReg1375_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1375_out;
SharedReg419_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg419_out;
SharedReg203_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg203_out;
SharedReg420_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg420_out;
SharedReg1049_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1049_out;
SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg210_out;
SharedReg1051_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1051_out;
SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg205_out;
SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg210_out;
SharedReg211_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg211_out;
SharedReg1648_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1648_out;
SharedReg1295_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1295_out;
SharedReg1059_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1059_out;
SharedReg1640_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1640_out;
SharedReg240_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg240_out;
SharedReg242_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg242_out;
SharedReg1594_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1594_out;
SharedReg218_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg218_out;
SharedReg1301_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1301_out;
SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg432_out;
SharedReg1379_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1379_out;
SharedReg1381_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1381_out;
SharedReg1601_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1601_out;
SharedReg1067_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1067_out;
   MUX_Product4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1633_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1389_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg396_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1373_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1374_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg183_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg427_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1028_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg220_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1380_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg189_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg403_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg404_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg434_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg439_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1383_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg184_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1032_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1566_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg426_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1375_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg419_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1628_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg203_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg420_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1049_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1051_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg210_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg211_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg438_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1648_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1295_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1059_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1640_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg240_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg242_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1594_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg218_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1301_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg432_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1071_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1379_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1381_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1601_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1067_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1576_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg193_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_6_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product4_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_7_impl_out,
                 X => Delay1No78_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1489_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1604_out;
SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1063_out;
SharedReg1600_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1600_out;
SharedReg1306_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1306_out;
SharedReg1631_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1548_out;
SharedReg1307_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1307_out;
SharedReg1524_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1635_out;
SharedReg219_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg219_out;
SharedReg1527_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1621_out;
SharedReg222_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg222_out;
SharedReg1517_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1537_out;
SharedReg1482_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1482_out;
SharedReg1086_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1086_out;
SharedReg1588_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1634_out;
SharedReg1298_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1298_out;
SharedReg1486_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1487_out;
SharedReg1091_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1091_out;
   MUX_Product4_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1489_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1630_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1548_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1307_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1524_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1641_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1635_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg219_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1527_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1528_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1498_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1499_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1490_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1500_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1501_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1502_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1591_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1503_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1504_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1593_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1556_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1506_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1507_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1603_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1508_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1509_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1510_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1560_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1511_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1512_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1513_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1514_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1565_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1621_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1604_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg222_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1517_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1518_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1519_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1520_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1610_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1532_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1582_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1534_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1535_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1521_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1522_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1585_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1536_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1523_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1537_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1482_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1086_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1588_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1634_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1600_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1298_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1486_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1487_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1091_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1306_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1631_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1495_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_7_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_7_impl_0_out,
                 Y => Delay1No78_out);

SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg1092_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1092_out;
SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg216_out;
SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1062_out;
SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1064_out;
SharedReg1601_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1601_out;
SharedReg1306_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg1633_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1633_out;
SharedReg1307_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1307_out;
SharedReg246_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg246_out;
SharedReg222_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg222_out;
SharedReg1628_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1628_out;
SharedReg221_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg221_out;
SharedReg1310_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1310_out;
SharedReg1311_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1311_out;
SharedReg1576_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1576_out;
SharedReg220_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg220_out;
SharedReg1072_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1072_out;
SharedReg426_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg426_out;
SharedReg1295_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1295_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg235_out;
SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg210_out;
SharedReg1296_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1296_out;
SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg210_out;
SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg236_out;
SharedReg1058_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1058_out;
SharedReg217_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg217_out;
SharedReg218_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg218_out;
SharedReg241_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg241_out;
SharedReg1302_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1302_out;
SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg216_out;
SharedReg433_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg433_out;
SharedReg434_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg434_out;
SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg213_out;
SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg243_out;
SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg213_out;
SharedReg1305_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1305_out;
SharedReg211_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg211_out;
SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1062_out;
SharedReg1566_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1566_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg235_out;
SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1297_out;
SharedReg448_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg448_out;
SharedReg228_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_48_cast <= SharedReg228_out;
SharedReg449_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg449_out;
SharedReg1078_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1078_out;
SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg261_out;
SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg261_out;
SharedReg1080_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1080_out;
SharedReg230_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg230_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_55_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg235_out;
SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg236_out;
SharedReg1648_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1648_out;
SharedReg1086_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1086_out;
SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1297_out;
SharedReg1640_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1640_out;
SharedReg266_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_62_cast <= SharedReg266_out;
SharedReg268_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg268_out;
SharedReg1594_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1594_out;
   MUX_Product4_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1092_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg222_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1628_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg221_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1310_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1311_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1576_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg220_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1072_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg426_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1295_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1296_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg210_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1058_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg217_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg218_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg241_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1302_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg216_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg433_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg434_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg243_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg213_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1305_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg211_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1062_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1566_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg448_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg228_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg449_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1078_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1601_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg261_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1080_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg230_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg235_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg236_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1648_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1086_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1297_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1640_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg266_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg268_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1594_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1633_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1307_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg246_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_7_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_7_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product4_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_8_impl_out,
                 X => Delay1No80_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1482_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1482_out;
SharedReg1457_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1457_out;
SharedReg1588_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1588_out;
SharedReg1634_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1634_out;
SharedReg1089_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1089_out;
SharedReg1486_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1486_out;
SharedReg1487_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1487_out;
SharedReg1462_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1462_out;
SharedReg1489_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1489_out;
SharedReg1630_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1630_out;
SharedReg1490_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1490_out;
SharedReg1603_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1603_out;
SharedReg1604_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1604_out;
SharedReg1093_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1093_out;
SharedReg1600_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1600_out;
SharedReg1097_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1097_out;
SharedReg1631_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1631_out;
SharedReg1495_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1548_out;
SharedReg1467_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1467_out;
SharedReg1524_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1524_out;
SharedReg1641_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1641_out;
SharedReg1635_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1635_out;
SharedReg271_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg271_out;
SharedReg1527_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1527_out;
SharedReg1528_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1528_out;
SharedReg1498_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1498_out;
SharedReg1499_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1499_out;
SharedReg1500_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1500_out;
SharedReg1501_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1501_out;
SharedReg1502_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1502_out;
SharedReg1591_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1591_out;
SharedReg1503_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1503_out;
SharedReg1504_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1504_out;
SharedReg1593_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1593_out;
SharedReg1556_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1556_out;
SharedReg1506_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1506_out;
SharedReg1507_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1507_out;
SharedReg1508_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1508_out;
SharedReg1509_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1509_out;
SharedReg1510_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1510_out;
SharedReg1560_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1560_out;
SharedReg1511_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1511_out;
SharedReg1512_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1512_out;
SharedReg1513_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1513_out;
SharedReg1514_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1514_out;
SharedReg1565_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1565_out;
SharedReg1621_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1621_out;
SharedReg274_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg274_out;
SharedReg1517_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1517_out;
SharedReg1518_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1518_out;
SharedReg1519_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1519_out;
SharedReg1520_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1520_out;
SharedReg1610_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1610_out;
SharedReg1532_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1532_out;
SharedReg1582_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1582_out;
SharedReg1534_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1534_out;
SharedReg1535_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1535_out;
SharedReg1521_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1521_out;
SharedReg1522_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1522_out;
SharedReg1585_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1585_out;
SharedReg1536_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1536_out;
SharedReg1523_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1523_out;
SharedReg1537_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1537_out;
   MUX_Product4_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1482_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1457_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1490_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1603_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1604_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1093_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1600_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1097_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1631_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1495_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1548_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1467_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1588_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1524_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1641_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1635_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg271_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1527_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1528_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1498_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1499_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1500_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1501_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1634_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1502_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1591_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1503_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1504_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1593_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1556_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1506_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1507_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1508_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1509_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1089_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1510_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1560_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1511_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1512_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1513_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1514_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1565_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1621_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg274_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1517_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1486_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1518_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1519_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1520_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1610_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1532_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1582_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1534_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1535_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1521_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1522_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1487_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1585_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1536_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1523_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1537_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1462_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1489_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1630_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_8_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_8_impl_0_out,
                 Y => Delay1No80_out);

SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg1648_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1648_out;
SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1457_out;
SharedReg1088_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1088_out;
SharedReg1640_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1640_out;
SharedReg461_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg461_out;
SharedReg463_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg463_out;
SharedReg1594_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1594_out;
SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg269_out;
SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1092_out;
SharedReg241_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg241_out;
SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1092_out;
SharedReg1303_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1303_out;
SharedReg1601_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1601_out;
SharedReg1306_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1306_out;
SharedReg1633_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1633_out;
SharedReg1098_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1098_out;
SharedReg467_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg467_out;
SharedReg274_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg274_out;
SharedReg1628_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1628_out;
SharedReg273_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg273_out;
SharedReg1470_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1470_out;
SharedReg1471_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1471_out;
SharedReg1576_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1576_out;
SharedReg272_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg272_out;
SharedReg1100_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1100_out;
SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg261_out;
SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1457_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg457_out;
SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg261_out;
SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg261_out;
SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1458_out;
SharedReg210_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg210_out;
SharedReg236_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg236_out;
SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1458_out;
SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg268_out;
SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg269_out;
SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg462_out;
SharedReg1093_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1093_out;
SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg462_out;
SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg268_out;
SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg269_out;
SharedReg213_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg213_out;
SharedReg464_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg464_out;
SharedReg264_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg264_out;
SharedReg1465_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1465_out;
SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg262_out;
SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1092_out;
SharedReg1566_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1566_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg457_out;
SharedReg1459_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1459_out;
SharedReg255_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_55_cast <= SharedReg255_out;
SharedReg478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg478_out;
SharedReg281_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg281_out;
SharedReg1476_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1476_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg457_out;
SharedReg1478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1478_out;
SharedReg282_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_62_cast <= SharedReg282_out;
SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_63_cast <= SharedReg261_out;
SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_64_cast <= SharedReg261_out;
   MUX_Product4_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1648_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg241_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1303_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1601_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1306_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1633_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1098_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg467_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg274_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1628_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg273_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1470_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1471_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1576_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg272_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1100_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1088_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg210_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg236_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1458_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1093_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg462_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1640_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg268_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg213_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg464_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg264_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1465_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg262_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1566_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg461_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1459_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg255_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg281_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1476_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg457_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg463_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1478_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg282_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg261_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1594_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg269_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1092_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_8_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_8_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product31_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_0_impl_out,
                 X => Delay1No82_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1535_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1571_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg1613_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1613_out;
SharedReg60_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg1537_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1540_out;
SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg297_out;
SharedReg295_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg295_out;
SharedReg1595_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1616_out;
SharedReg861_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg861_out;
SharedReg1492_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1494_out;
SharedReg301_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg301_out;
SharedReg1496_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1578_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg36_out;
SharedReg1400_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1400_out;
SharedReg1636_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1552_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg36_out;
SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1401_out;
SharedReg1554_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1554_out;
SharedReg291_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg291_out;
SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1401_out;
SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg297_out;
SharedReg1638_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1508_out;
SharedReg296_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg296_out;
SharedReg1639_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1562_out;
SharedReg39_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg39_out;
SharedReg1564_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1516_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg36_out;
SharedReg1569_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1625_out;
SharedReg58_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg58_out;
SharedReg1533_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1583_out;
   MUX_Product31_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1535_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1571_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1485_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1651_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1540_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg295_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1595_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1632_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1543_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1616_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg861_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1492_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1600_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1493_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1494_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg301_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1496_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1497_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1574_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1615_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1525_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1613_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1526_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1527_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1578_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1400_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1636_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1552_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1554_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg60_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg291_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1401_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg297_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1638_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1557_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1508_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg296_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1639_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1605_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1561_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1562_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg39_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1564_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1515_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1531_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1516_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1569_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1570_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1537_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1625_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg58_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1533_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1583_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1650_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1483_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1646_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_0_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_0_impl_0_out,
                 Y => Delay1No82_out);

SharedReg874_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg874_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg1572_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1572_out;
SharedReg854_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg854_out;
SharedReg1586_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1573_out;
SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg853_out;
SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg853_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg1401_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1401_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg857_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg857_out;
SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg41_out;
SharedReg1541_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1542_out;
SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg859_out;
SharedReg1406_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1406_out;
SharedReg295_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg295_out;
SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg859_out;
SharedReg1617_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1617_out;
SharedReg45_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg45_out;
SharedReg861_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg861_out;
SharedReg300_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg300_out;
SharedReg302_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg302_out;
SharedReg1547_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1547_out;
SharedReg305_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg305_out;
SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg47_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg47_out;
SharedReg1413_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1413_out;
SharedReg303_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg303_out;
SharedReg1414_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1414_out;
SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg49_out;
SharedReg866_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg866_out;
SharedReg1550_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1551_out;
SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg853_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg36_out;
SharedReg1553_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1597_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg36_out;
SharedReg1555_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1556_out;
SharedReg1408_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1408_out;
SharedReg296_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg296_out;
SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg859_out;
SharedReg1559_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1559_out;
SharedReg860_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg860_out;
SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg859_out;
SharedReg39_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg39_out;
SharedReg298_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg298_out;
SharedReg1563_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1563_out;
SharedReg1410_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1410_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg37_out;
SharedReg1420_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1420_out;
SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg48_out;
SharedReg1567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1568_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg36_out;
SharedReg855_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg855_out;
SharedReg1581_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1581_out;
SharedReg1421_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1421_out;
SharedReg59_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg59_out;
   MUX_Product31_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg874_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg857_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1541_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1542_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1406_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg295_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1617_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1572_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg45_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg861_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg300_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg302_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1547_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg305_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg47_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1413_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg303_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg854_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1414_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg866_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1550_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1551_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1553_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1597_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1586_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1555_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1599_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1556_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1408_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg296_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1559_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg860_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg859_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg39_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg298_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1563_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1410_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1420_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg48_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg855_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1581_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1421_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg59_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg853_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1401_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_0_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_0_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product31_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_1_impl_out,
                 X => Delay1No84_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast);

SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg1569_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1625_out;
SharedReg311_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg311_out;
SharedReg1533_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1571_out;
SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg66_out;
SharedReg1613_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1613_out;
SharedReg89_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg66_out;
SharedReg1537_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1540_out;
SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg324_out;
SharedReg322_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg322_out;
SharedReg1595_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1616_out;
SharedReg890_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg890_out;
SharedReg1492_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1494_out;
SharedReg328_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg328_out;
SharedReg1496_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1578_out;
SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg66_out;
SharedReg1347_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1347_out;
SharedReg1636_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1552_out;
SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg66_out;
SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1348_out;
SharedReg1554_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1554_out;
SharedReg318_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg318_out;
SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1348_out;
SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg324_out;
SharedReg1638_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1508_out;
SharedReg323_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg323_out;
SharedReg1639_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1562_out;
SharedReg293_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg293_out;
SharedReg1564_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1516_out;
SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg290_out;
   MUX_Product31_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1569_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1613_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1537_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1650_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1483_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1646_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1485_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1651_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1540_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1570_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg322_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1595_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1632_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1543_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1616_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg890_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1492_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1600_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1493_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1625_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1494_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg328_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1496_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1497_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1574_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1615_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1525_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1526_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1527_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1578_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg311_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1347_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1636_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1552_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1554_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg318_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1348_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg324_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1533_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1638_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1557_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1508_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg323_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1639_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1605_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1561_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1562_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg293_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1564_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1583_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1515_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1531_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1516_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg290_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1535_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1571_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_1_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_0_out,
                 Y => Delay1No84_out);

SharedReg1568_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1568_out;
SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg1402_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1402_out;
SharedReg1581_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1581_out;
SharedReg1366_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1366_out;
SharedReg88_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg902_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg902_out;
SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg66_out;
SharedReg1572_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1572_out;
SharedReg883_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg883_out;
SharedReg1586_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1573_out;
SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg882_out;
SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg882_out;
SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg66_out;
SharedReg1348_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1348_out;
SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg67_out;
SharedReg886_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg886_out;
SharedReg71_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg71_out;
SharedReg1541_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1542_out;
SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg888_out;
SharedReg1353_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1353_out;
SharedReg322_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg322_out;
SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg888_out;
SharedReg1617_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1617_out;
SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg75_out;
SharedReg890_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg890_out;
SharedReg327_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg327_out;
SharedReg329_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg329_out;
SharedReg1547_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1547_out;
SharedReg332_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg332_out;
SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg78_out;
SharedReg77_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg77_out;
SharedReg1360_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1360_out;
SharedReg330_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg330_out;
SharedReg1361_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1361_out;
SharedReg79_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg79_out;
SharedReg895_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg895_out;
SharedReg1550_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1551_out;
SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg882_out;
SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg66_out;
SharedReg1553_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1597_out;
SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg66_out;
SharedReg1555_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1556_out;
SharedReg1355_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1355_out;
SharedReg323_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg323_out;
SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg888_out;
SharedReg1559_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1559_out;
SharedReg889_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg889_out;
SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg888_out;
SharedReg69_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg69_out;
SharedReg325_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg325_out;
SharedReg1563_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1563_out;
SharedReg1357_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1357_out;
SharedReg291_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg291_out;
SharedReg1365_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1365_out;
SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg78_out;
SharedReg1567_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1567_out;
   MUX_Product31_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1568_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg883_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1586_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1573_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1348_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg886_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg71_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg290_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1541_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1542_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1353_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg322_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1617_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg890_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg327_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1402_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg329_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1547_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg332_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg77_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1360_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg330_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1361_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg79_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg895_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1581_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1550_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1551_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg882_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1553_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1555_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1556_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1366_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1355_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg323_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1559_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg889_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg888_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg69_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg325_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1563_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1357_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg291_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1365_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg78_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1567_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg902_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg66_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1572_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_1_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product31_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_2_impl_out,
                 X => Delay1No86_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1562_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1562_out;
SharedReg69_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg1564_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1516_out;
SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg317_out;
SharedReg1569_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1625_out;
SharedReg336_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg336_out;
SharedReg1533_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1571_out;
SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg1613_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1613_out;
SharedReg117_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg117_out;
SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg95_out;
SharedReg1537_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1540_out;
SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg350_out;
SharedReg348_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg348_out;
SharedReg1595_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1616_out;
SharedReg918_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg918_out;
SharedReg1492_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1494_out;
SharedReg354_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg354_out;
SharedReg1496_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1578_out;
SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg95_out;
SharedReg1428_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1428_out;
SharedReg1636_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1552_out;
SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg95_out;
SharedReg1429_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1429_out;
SharedReg1554_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1554_out;
SharedReg344_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg344_out;
SharedReg911_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg911_out;
SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg350_out;
SharedReg1638_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1508_out;
SharedReg101_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg101_out;
SharedReg1639_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1561_out;
   MUX_Product31_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1562_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg336_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1533_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1583_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1535_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1571_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1613_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg117_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1564_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1537_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1650_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1483_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1646_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1485_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1651_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1540_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg348_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1595_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1515_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1632_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1543_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1616_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg918_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1492_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1600_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1493_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1494_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg354_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1496_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1531_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1497_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1574_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1615_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1525_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1526_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1527_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1578_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1428_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1636_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1516_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1552_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg95_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1429_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1554_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg344_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg911_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg350_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1638_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1557_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1508_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg101_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1639_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1605_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1561_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg317_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1569_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1570_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_2_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_2_impl_0_out,
                 Y => Delay1No86_out);

SharedReg103_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg1563_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1563_out;
SharedReg920_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg67_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg67_out;
SharedReg1446_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1446_out;
SharedReg330_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg330_out;
SharedReg1567_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1568_out;
SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg1349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1349_out;
SharedReg1581_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1581_out;
SharedReg1447_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1447_out;
SharedReg116_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg116_out;
SharedReg930_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg930_out;
SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg95_out;
SharedReg1572_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1572_out;
SharedReg911_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg911_out;
SharedReg1586_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1573_out;
SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg910_out;
SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg910_out;
SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg95_out;
SharedReg1429_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1429_out;
SharedReg96_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg96_out;
SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg914_out;
SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg100_out;
SharedReg1541_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1542_out;
SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg916_out;
SharedReg1434_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1434_out;
SharedReg348_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg348_out;
SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg916_out;
SharedReg1617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1617_out;
SharedReg104_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg104_out;
SharedReg918_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg918_out;
SharedReg353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg353_out;
SharedReg355_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg355_out;
SharedReg1547_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1547_out;
SharedReg358_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg358_out;
SharedReg107_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg107_out;
SharedReg106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg106_out;
SharedReg1441_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1441_out;
SharedReg356_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg356_out;
SharedReg1442_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1442_out;
SharedReg108_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg108_out;
SharedReg923_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg923_out;
SharedReg1550_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1551_out;
SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg910_out;
SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg95_out;
SharedReg1553_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1597_out;
SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg95_out;
SharedReg1555_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1556_out;
SharedReg1436_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1436_out;
SharedReg349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg349_out;
SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1353_out;
SharedReg1559_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1559_out;
SharedReg1354_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1354_out;
SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1353_out;
SharedReg320_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg320_out;
   MUX_Product31_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1563_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1581_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1447_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg116_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg930_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1572_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg911_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1586_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1573_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1429_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg96_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1541_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1542_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg67_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1434_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg348_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg916_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg104_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg918_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg355_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1547_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg358_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1446_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg107_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1441_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg356_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1442_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg108_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg923_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1550_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1551_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg910_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg330_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1553_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1597_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1555_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1599_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1556_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1436_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg349_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1567_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1559_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1354_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1353_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg320_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1568_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_2_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_2_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product31_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_3_impl_out,
                 X => Delay1No88_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1638_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1508_out;
SharedReg349_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
SharedReg1639_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1562_out;
SharedReg98_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg98_out;
SharedReg1564_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1516_out;
SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg343_out;
SharedReg1569_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1625_out;
SharedReg362_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg362_out;
SharedReg1533_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1571_out;
SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg124_out;
SharedReg1613_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1613_out;
SharedReg146_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg146_out;
SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg124_out;
SharedReg1537_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1540_out;
SharedReg375_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg375_out;
SharedReg373_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg373_out;
SharedReg1595_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1616_out;
SharedReg948_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg948_out;
SharedReg1492_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1494_out;
SharedReg379_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg379_out;
SharedReg1496_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1578_out;
SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg343_out;
SharedReg940_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg940_out;
SharedReg1636_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1552_out;
SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg343_out;
SharedReg941_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg941_out;
SharedReg1554_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1554_out;
SharedReg125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg125_out;
SharedReg1429_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1429_out;
SharedReg131_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg131_out;
   MUX_Product31_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1638_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1557_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1515_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1531_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1516_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1569_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1570_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1625_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg362_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1533_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1508_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1583_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1535_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1571_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1613_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg146_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1537_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1650_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1483_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1646_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1485_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1651_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1540_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg375_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg373_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1595_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1632_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1543_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1616_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1639_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg948_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1492_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1600_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1493_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1494_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg379_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1496_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1497_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1574_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1615_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1605_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1525_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1526_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1527_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1578_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg940_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1636_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1552_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg343_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg941_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1561_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1554_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1429_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg131_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1562_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg98_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1564_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_3_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_0_out,
                 Y => Delay1No88_out);

SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg948_out;
SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg1559_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1559_out;
SharedReg917_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg916_out;
SharedReg98_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg98_out;
SharedReg351_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg351_out;
SharedReg1563_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1563_out;
SharedReg1438_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1438_out;
SharedReg96_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg1339_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1339_out;
SharedReg107_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg107_out;
SharedReg1567_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1568_out;
SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg343_out;
SharedReg1430_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1430_out;
SharedReg1581_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1581_out;
SharedReg1340_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1340_out;
SharedReg145_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg145_out;
SharedReg960_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg960_out;
SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg124_out;
SharedReg1572_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1572_out;
SharedReg941_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg941_out;
SharedReg1586_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1573_out;
SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg940_out;
SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg940_out;
SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg124_out;
SharedReg1322_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1322_out;
SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg125_out;
SharedReg944_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg944_out;
SharedReg129_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg129_out;
SharedReg1541_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1542_out;
SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg946_out;
SharedReg1327_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1327_out;
SharedReg373_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg373_out;
SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg946_out;
SharedReg1617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1617_out;
SharedReg133_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg133_out;
SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg948_out;
SharedReg378_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg378_out;
SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg135_out;
SharedReg1547_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1547_out;
SharedReg383_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg383_out;
SharedReg136_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg136_out;
SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg135_out;
SharedReg1334_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1334_out;
SharedReg381_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg381_out;
SharedReg1335_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1335_out;
SharedReg137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg137_out;
SharedReg953_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg953_out;
SharedReg1550_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1551_out;
SharedReg1428_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1428_out;
SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg343_out;
SharedReg1553_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1597_out;
SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg343_out;
SharedReg1555_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1556_out;
   MUX_Product31_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1339_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg107_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1567_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1568_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1430_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1581_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1340_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg145_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg960_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1572_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg941_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1586_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1573_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg940_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg124_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1559_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1322_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg944_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg129_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1541_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1542_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1327_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg373_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg946_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg917_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg133_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg948_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg378_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1547_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg383_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg136_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg135_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1334_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg381_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1335_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg953_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1550_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1551_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1428_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1553_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1597_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg98_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg343_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1555_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1599_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1556_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg351_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1563_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1438_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_3_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product31_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_4_impl_out,
                 X => Delay1No90_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1552_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1552_out;
SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg124_out;
SharedReg1322_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1322_out;
SharedReg1554_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1554_out;
SharedReg369_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg369_out;
SharedReg941_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg941_out;
SharedReg375_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg375_out;
SharedReg1638_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1508_out;
SharedReg130_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg130_out;
SharedReg1639_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1562_out;
SharedReg127_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg127_out;
SharedReg1564_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1516_out;
SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg368_out;
SharedReg1569_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1625_out;
SharedReg388_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg388_out;
SharedReg1533_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1571_out;
SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg154_out;
SharedReg1613_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1613_out;
SharedReg390_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg390_out;
SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg154_out;
SharedReg1537_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1540_out;
SharedReg403_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg403_out;
SharedReg401_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg401_out;
SharedReg1595_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1616_out;
SharedReg976_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg976_out;
SharedReg1492_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1494_out;
SharedReg407_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg407_out;
SharedReg1496_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1578_out;
SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg124_out;
SharedReg1321_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1321_out;
SharedReg1636_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1636_out;
   MUX_Product31_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1552_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg130_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1639_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1605_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1561_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1562_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg127_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1564_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1515_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1531_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1322_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg368_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1569_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1570_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1625_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg388_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1533_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1583_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1535_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1571_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1554_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1613_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg390_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg154_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1537_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1650_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1483_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1646_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1485_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1651_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg369_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1540_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg403_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg401_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1595_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1632_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1543_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1616_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg976_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1492_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1600_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg941_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1493_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1494_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg407_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1496_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1497_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1574_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1615_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1525_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1526_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1527_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg375_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1578_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg124_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1321_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1636_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1638_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1557_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1508_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_4_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_0_out,
                 Y => Delay1No90_out);

SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg1553_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1597_out;
SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg1555_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1556_out;
SharedReg1329_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1329_out;
SharedReg374_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg374_out;
SharedReg1434_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1434_out;
SharedReg1559_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1559_out;
SharedReg1435_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1435_out;
SharedReg946_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg946_out;
SharedReg127_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
SharedReg376_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg376_out;
SharedReg1563_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1563_out;
SharedReg1331_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1331_out;
SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg125_out;
SharedReg1019_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1019_out;
SharedReg136_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg136_out;
SharedReg1567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1568_out;
SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg368_out;
SharedReg1323_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1323_out;
SharedReg1581_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1581_out;
SharedReg988_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg988_out;
SharedReg389_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg389_out;
SharedReg1341_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1341_out;
SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg154_out;
SharedReg1572_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1572_out;
SharedReg969_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg969_out;
SharedReg1586_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1573_out;
SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg968_out;
SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg968_out;
SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg154_out;
SharedReg999_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg999_out;
SharedReg155_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg155_out;
SharedReg972_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg972_out;
SharedReg159_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg159_out;
SharedReg1541_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1542_out;
SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg974_out;
SharedReg1004_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1004_out;
SharedReg401_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg401_out;
SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg974_out;
SharedReg1617_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1617_out;
SharedReg164_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg164_out;
SharedReg976_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg976_out;
SharedReg406_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg406_out;
SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg166_out;
SharedReg1547_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1547_out;
SharedReg411_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg411_out;
SharedReg167_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg167_out;
SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg166_out;
SharedReg1011_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1011_out;
SharedReg409_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg409_out;
SharedReg1012_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1012_out;
SharedReg168_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg168_out;
SharedReg981_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg981_out;
SharedReg1550_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1551_out;
SharedReg940_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg940_out;
   MUX_Product31_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1553_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1559_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1435_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg946_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg376_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1563_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1331_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1019_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg136_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1597_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1568_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg368_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1323_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1581_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg988_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg389_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1341_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg124_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1572_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg969_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1586_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1573_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg968_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg154_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg999_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg155_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg972_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1555_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg159_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1541_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1542_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1004_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg401_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg974_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1617_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg164_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg976_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1599_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg406_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1547_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg411_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg167_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg166_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1011_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg409_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1012_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg168_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1556_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg981_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1550_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1551_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg940_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1329_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg374_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1434_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_4_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product31_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_5_impl_out,
                 X => Delay1No92_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1525_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1578_out;
SharedReg368_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg998_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1636_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1552_out;
SharedReg154_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg154_out;
SharedReg999_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg999_out;
SharedReg1554_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1554_out;
SharedReg397_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg397_out;
SharedReg969_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg969_out;
SharedReg403_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg403_out;
SharedReg1638_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1508_out;
SharedReg160_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg160_out;
SharedReg1639_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1562_out;
SharedReg157_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg157_out;
SharedReg1564_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1516_out;
SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg396_out;
SharedReg1569_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1625_out;
SharedReg176_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg176_out;
SharedReg1533_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1571_out;
SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg183_out;
SharedReg1613_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1613_out;
SharedReg178_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg178_out;
SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg183_out;
SharedReg1537_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1540_out;
SharedReg433_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg433_out;
SharedReg431_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg431_out;
SharedReg1595_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1616_out;
SharedReg1034_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1034_out;
SharedReg1492_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1494_out;
SharedReg437_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg437_out;
SharedReg1496_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1615_out;
   MUX_Product31_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1525_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1526_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1554_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg397_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg969_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg403_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1638_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1557_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1508_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg160_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1639_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1605_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1527_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1561_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1562_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg157_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1564_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1515_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1531_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1516_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg396_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1569_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1578_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1570_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1625_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg176_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1533_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1583_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1535_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1571_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1613_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg178_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg368_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg183_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1537_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1650_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1483_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1646_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1485_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1651_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1540_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg433_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg431_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg998_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1595_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1632_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1543_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1616_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1034_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1492_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1600_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1493_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1494_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg437_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1636_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1496_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1497_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1574_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1615_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1552_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg154_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg999_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_5_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_5_impl_0_out,
                 Y => Delay1No92_out);

SharedReg439_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg439_out;
SharedReg1387_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1387_out;
SharedReg197_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg197_out;
SharedReg1040_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1040_out;
SharedReg1550_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1551_out;
SharedReg968_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg968_out;
SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg154_out;
SharedReg1553_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1597_out;
SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg154_out;
SharedReg1555_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1556_out;
SharedReg1006_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1006_out;
SharedReg402_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg402_out;
SharedReg1327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1327_out;
SharedReg1559_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1559_out;
SharedReg1328_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1328_out;
SharedReg974_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg974_out;
SharedReg157_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg157_out;
SharedReg404_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg404_out;
SharedReg1563_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1563_out;
SharedReg1008_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1008_out;
SharedReg155_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg155_out;
SharedReg1047_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1047_out;
SharedReg167_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg167_out;
SharedReg1567_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1568_out;
SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg396_out;
SharedReg1000_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1000_out;
SharedReg1581_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1581_out;
SharedReg1020_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1020_out;
SharedReg177_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg177_out;
SharedReg989_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg989_out;
SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg183_out;
SharedReg1572_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1572_out;
SharedReg1028_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1028_out;
SharedReg1586_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1573_out;
SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1027_out;
SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1027_out;
SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg183_out;
SharedReg1374_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1374_out;
SharedReg184_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg184_out;
SharedReg1031_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1031_out;
SharedReg188_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg188_out;
SharedReg1541_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1542_out;
SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1032_out;
SharedReg1379_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1379_out;
SharedReg431_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg431_out;
SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1032_out;
SharedReg1617_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1617_out;
SharedReg192_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg192_out;
SharedReg1034_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1034_out;
SharedReg436_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg436_out;
SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg194_out;
SharedReg1547_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1547_out;
SharedReg441_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg441_out;
SharedReg195_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg195_out;
SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg194_out;
SharedReg1386_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1386_out;
   MUX_Product31_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg439_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1387_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1555_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1599_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1556_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1006_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg402_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1559_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1328_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg974_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg197_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg157_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg404_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1563_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1008_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg155_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1047_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg167_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1567_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1568_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1040_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg396_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1000_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1581_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1020_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg177_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg989_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1572_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1028_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1586_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1550_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1573_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1027_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg183_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1374_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg184_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1031_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg188_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1541_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1542_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1551_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1379_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg431_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1032_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1617_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg192_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1034_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg436_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1547_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg968_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg441_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg195_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg194_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1386_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg154_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1553_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1597_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_5_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_5_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product31_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_6_impl_out,
                 X => Delay1No94_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1493_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1494_out;
SharedReg220_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg1496_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1578_out;
SharedReg396_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg396_out;
SharedReg1373_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1373_out;
SharedReg1636_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1552_out;
SharedReg183_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg183_out;
SharedReg1374_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1374_out;
SharedReg1554_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1554_out;
SharedReg427_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg427_out;
SharedReg1028_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1028_out;
SharedReg433_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg433_out;
SharedReg1638_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1508_out;
SharedReg189_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg189_out;
SharedReg1639_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1562_out;
SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg186_out;
SharedReg1564_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1516_out;
SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg426_out;
SharedReg1569_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1625_out;
SharedReg419_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg419_out;
SharedReg1533_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1571_out;
SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg210_out;
SharedReg1613_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1613_out;
SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg205_out;
SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg210_out;
SharedReg1537_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1540_out;
SharedReg242_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg242_out;
SharedReg240_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg240_out;
SharedReg1595_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1616_out;
SharedReg1381_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1381_out;
SharedReg1492_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1600_out;
   MUX_Product31_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1493_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1494_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1578_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg396_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1373_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1636_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1552_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg183_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1374_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1554_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg427_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1028_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg220_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg433_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1638_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1557_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1508_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg189_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1639_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1605_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1561_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1562_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1496_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1564_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1515_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1531_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1516_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg426_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1569_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1570_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1625_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg419_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1497_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1533_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1583_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1535_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1571_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1613_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg210_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1537_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1650_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1574_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1483_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1646_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1485_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1651_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1540_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg242_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg240_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1595_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1632_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1543_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1615_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1616_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1381_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1492_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1600_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1525_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1526_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1527_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_6_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_6_impl_0_out,
                 Y => Delay1No94_out);

SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg219_out;
SharedReg221_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg1547_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1547_out;
SharedReg250_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg250_out;
SharedReg439_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg439_out;
SharedReg438_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
SharedReg1069_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1069_out;
SharedReg222_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg222_out;
SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1070_out;
SharedReg441_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg441_out;
SharedReg1389_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1389_out;
SharedReg1550_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1551_out;
SharedReg1027_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1027_out;
SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg183_out;
SharedReg1553_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1597_out;
SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg183_out;
SharedReg1555_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1556_out;
SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1381_out;
SharedReg432_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg432_out;
SharedReg1004_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1004_out;
SharedReg1559_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1559_out;
SharedReg1005_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1005_out;
SharedReg1032_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1032_out;
SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg186_out;
SharedReg434_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg434_out;
SharedReg1563_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1563_out;
SharedReg1383_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1383_out;
SharedReg184_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg184_out;
SharedReg1393_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1393_out;
SharedReg195_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg195_out;
SharedReg1567_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1568_out;
SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg426_out;
SharedReg1375_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1375_out;
SharedReg1581_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1581_out;
SharedReg1048_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1048_out;
SharedReg420_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg420_out;
SharedReg1021_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1021_out;
SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg210_out;
SharedReg1572_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1572_out;
SharedReg1058_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1058_out;
SharedReg1586_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1573_out;
SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1057_out;
SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1057_out;
SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg210_out;
SharedReg1296_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1296_out;
SharedReg211_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg211_out;
SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1061_out;
SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg215_out;
SharedReg1541_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1542_out;
SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1062_out;
SharedReg1301_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1301_out;
SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg215_out;
SharedReg1379_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1379_out;
SharedReg1617_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1617_out;
SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg219_out;
SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1381_out;
   MUX_Product31_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1389_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1550_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1551_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1027_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1553_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1597_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg183_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1555_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1599_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1547_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1556_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg432_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1004_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1559_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1005_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1032_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg434_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1563_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg250_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1383_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg184_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1393_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg195_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1567_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1568_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg426_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1375_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1581_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg439_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1048_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg420_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1021_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1572_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1058_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1586_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1573_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1057_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg438_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg210_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1296_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg211_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1541_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1542_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1301_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg215_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1069_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1379_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1617_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg219_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1381_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg222_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg441_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_6_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_6_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product31_7_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product31_7_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product31_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_7_impl_out,
                 X => Delay1No96_out_to_Product31_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product31_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1595_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1616_out;
SharedReg1064_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1064_out;
SharedReg1492_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1494_out;
SharedReg246_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg246_out;
SharedReg1496_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1578_out;
SharedReg426_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg426_out;
SharedReg1295_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1295_out;
SharedReg1636_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1552_out;
SharedReg210_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg210_out;
SharedReg1296_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1296_out;
SharedReg1554_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1554_out;
SharedReg236_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg236_out;
SharedReg1058_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1058_out;
SharedReg242_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg242_out;
SharedReg1638_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1508_out;
SharedReg216_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg216_out;
SharedReg1639_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1562_out;
SharedReg213_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg213_out;
SharedReg1564_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1516_out;
SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg235_out;
SharedReg1569_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1625_out;
SharedReg448_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg448_out;
SharedReg1533_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1571_out;
SharedReg261_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg261_out;
SharedReg1613_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1613_out;
SharedReg230_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg230_out;
SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg235_out;
SharedReg1537_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1537_out;
SharedReg1650_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1540_out;
SharedReg268_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg268_out;
SharedReg266_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg266_out;
   MUX_Product31_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1595_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1632_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1496_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1497_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1574_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1615_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1525_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1526_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1527_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1578_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg426_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1295_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1543_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1636_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1552_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg210_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1296_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1554_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg236_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1058_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg242_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1638_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1557_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1616_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1508_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg216_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1639_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1605_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1561_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1562_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg213_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1564_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1515_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1531_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1064_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1516_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1569_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1570_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1625_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg448_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1533_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1583_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1535_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1492_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1571_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg261_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1613_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg230_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg235_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1537_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1650_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1483_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1646_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1485_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1600_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1651_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1540_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg268_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg266_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1493_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1494_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg246_out_to_MUX_Product31_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_7_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_7_impl_0_out,
                 Y => Delay1No96_out);

SharedReg1301_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1301_out;
SharedReg1092_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1092_out;
SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg240_out;
SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1062_out;
SharedReg1617_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1617_out;
SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg245_out;
SharedReg1064_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1064_out;
SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg245_out;
SharedReg247_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg247_out;
SharedReg1547_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1547_out;
SharedReg276_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg276_out;
SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg222_out;
SharedReg221_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg221_out;
SharedReg1308_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1308_out;
SharedReg248_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg248_out;
SharedReg1309_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1309_out;
SharedReg223_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg223_out;
SharedReg1072_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1072_out;
SharedReg1550_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1551_out;
SharedReg1057_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1057_out;
SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg1553_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1597_out;
SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg210_out;
SharedReg1555_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1556_out;
SharedReg1303_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1303_out;
SharedReg241_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg241_out;
SharedReg1379_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1379_out;
SharedReg1559_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1559_out;
SharedReg1380_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1380_out;
SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1062_out;
SharedReg213_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg213_out;
SharedReg243_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg243_out;
SharedReg1563_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1563_out;
SharedReg1305_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1305_out;
SharedReg211_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg211_out;
SharedReg1313_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1313_out;
SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg222_out;
SharedReg1567_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1568_out;
SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg235_out;
SharedReg1297_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1297_out;
SharedReg1581_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1581_out;
SharedReg1077_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1077_out;
SharedReg449_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg449_out;
SharedReg1394_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1394_out;
SharedReg261_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg261_out;
SharedReg1572_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1572_out;
SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1087_out;
SharedReg1586_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1573_out;
SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1295_out;
SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1295_out;
SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg235_out;
SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1087_out;
SharedReg236_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_60_cast <= SharedReg236_out;
SharedReg1299_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1299_out;
SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_62_cast <= SharedReg240_out;
SharedReg1541_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1542_out;
   MUX_Product31_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1301_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1092_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg221_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1308_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg248_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1309_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg223_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1072_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1550_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1551_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1057_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1553_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1597_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg210_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1555_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1599_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1556_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1303_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg241_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1379_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1559_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1380_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1062_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg213_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg243_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1563_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1305_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg211_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1313_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1617_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg222_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1567_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1568_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1297_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1581_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1077_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg449_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1394_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg261_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1572_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1586_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1573_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1295_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg235_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1087_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg236_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1064_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1299_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg240_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1541_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1542_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg245_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg247_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1547_out_to_MUX_Product31_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_7_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_7_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product31_8_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product31_8_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product31_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_8_impl_out,
                 X => Delay1No98_out_to_Product31_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product31_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1650_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1650_out;
SharedReg1483_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1483_out;
SharedReg1646_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1646_out;
SharedReg1485_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1485_out;
SharedReg1651_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1540_out;
SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg463_out;
SharedReg461_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg461_out;
SharedReg1595_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1595_out;
SharedReg1632_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1632_out;
SharedReg1543_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1543_out;
SharedReg1616_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1616_out;
SharedReg1303_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1303_out;
SharedReg1492_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1492_out;
SharedReg1600_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1600_out;
SharedReg1493_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1493_out;
SharedReg1494_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1494_out;
SharedReg467_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg467_out;
SharedReg1496_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1496_out;
SharedReg1497_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1497_out;
SharedReg1574_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1574_out;
SharedReg1615_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1615_out;
SharedReg1525_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1525_out;
SharedReg1526_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1526_out;
SharedReg1527_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1527_out;
SharedReg1578_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1578_out;
SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg261_out;
SharedReg1457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1457_out;
SharedReg1636_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1636_out;
SharedReg1552_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1552_out;
SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg261_out;
SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1458_out;
SharedReg1554_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1554_out;
SharedReg236_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg236_out;
SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1458_out;
SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg463_out;
SharedReg1638_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1638_out;
SharedReg1557_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1557_out;
SharedReg1508_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1508_out;
SharedReg462_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg462_out;
SharedReg1639_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1639_out;
SharedReg1605_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1605_out;
SharedReg1561_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1561_out;
SharedReg1562_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1562_out;
SharedReg264_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg264_out;
SharedReg1564_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1564_out;
SharedReg1515_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1515_out;
SharedReg1531_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1531_out;
SharedReg1516_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1516_out;
SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg457_out;
SharedReg1569_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1569_out;
SharedReg1570_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1570_out;
SharedReg1625_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1625_out;
SharedReg255_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg255_out;
SharedReg1533_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1533_out;
SharedReg1583_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1583_out;
SharedReg1535_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1535_out;
SharedReg1571_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1571_out;
SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg457_out;
SharedReg1613_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1613_out;
SharedReg282_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_62_cast <= SharedReg282_out;
SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_63_cast <= SharedReg261_out;
SharedReg1537_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1537_out;
   MUX_Product31_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1650_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1483_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1543_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1616_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1303_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1492_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1600_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1493_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1494_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg467_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1496_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1497_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1646_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1574_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1615_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1525_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1526_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1527_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1578_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1636_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1552_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1485_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1554_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg236_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1458_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1638_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1557_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1508_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg462_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1651_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1639_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1605_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1561_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1562_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg264_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1564_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1515_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1531_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1516_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1540_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1569_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1570_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1625_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg255_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1533_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1583_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1535_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1571_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg457_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg463_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1613_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg282_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg261_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1537_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg461_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1595_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1632_out_to_MUX_Product31_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_8_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_8_impl_0_out,
                 Y => Delay1No98_out);

SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1086_out;
SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg261_out;
SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1458_out;
SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg1090_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1090_out;
SharedReg266_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg266_out;
SharedReg1541_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1541_out;
SharedReg1542_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1542_out;
SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1092_out;
SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1092_out;
SharedReg461_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg461_out;
SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1092_out;
SharedReg1617_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1617_out;
SharedReg245_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg245_out;
SharedReg1094_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1094_out;
SharedReg466_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg466_out;
SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg273_out;
SharedReg1547_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1547_out;
SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg276_out;
SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg274_out;
SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg273_out;
SharedReg1468_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1468_out;
SharedReg469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg469_out;
SharedReg1469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1469_out;
SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg276_out;
SharedReg1100_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1100_out;
SharedReg1550_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1550_out;
SharedReg1551_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1551_out;
SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1086_out;
SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg261_out;
SharedReg1553_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1553_out;
SharedReg1597_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1597_out;
SharedReg210_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg210_out;
SharedReg1555_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1555_out;
SharedReg1599_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1599_out;
SharedReg1556_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1556_out;
SharedReg1463_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1463_out;
SharedReg462_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg462_out;
SharedReg1301_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1301_out;
SharedReg1559_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1559_out;
SharedReg1093_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1093_out;
SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1092_out;
SharedReg213_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg213_out;
SharedReg464_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg464_out;
SharedReg1563_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1563_out;
SharedReg1465_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1465_out;
SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg262_out;
SharedReg1475_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1475_out;
SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg274_out;
SharedReg1567_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1567_out;
SharedReg1568_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1568_out;
SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg457_out;
SharedReg1459_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1459_out;
SharedReg1581_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1581_out;
SharedReg1106_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1106_out;
SharedReg281_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg281_out;
SharedReg1107_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1107_out;
SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg457_out;
SharedReg1572_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1572_out;
SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1458_out;
SharedReg1586_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1586_out;
SharedReg1573_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1573_out;
SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1086_out;
   MUX_Product31_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg461_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1617_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg245_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1094_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg466_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1547_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg273_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1468_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1469_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg276_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1100_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1550_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1551_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg261_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1553_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1597_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg210_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1555_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1599_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1556_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1463_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg462_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1301_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1559_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1090_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1093_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg213_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg464_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1563_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1465_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg262_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1475_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg274_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1567_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg266_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1568_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1459_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1581_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1106_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg281_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1107_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg457_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1572_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1541_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1458_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1586_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1573_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1086_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1542_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1092_out_to_MUX_Product31_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_8_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_8_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No100_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg484_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg488_out;
SharedReg496_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg496_out;
SharedReg864_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg864_out;
SharedReg1129_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1129_out;
SharedReg688_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg688_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg673_out;
SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg677_out;
SharedReg684_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg684_out;
SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg490_out;
SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1116_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg484_out;
SharedReg1115_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1115_out;
SharedReg872_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg872_out;
SharedReg1403_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1403_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg485_out;
SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg295_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg484_out;
SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg490_out;
SharedReg1130_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1130_out;
SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg677_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg673_out;
SharedReg853_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg853_out;
SharedReg1131_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1131_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg485_out;
SharedReg290_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg290_out;
SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg302_out;
SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg855_out;
SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg487_out;
SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg52_out;
SharedReg676_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg676_out;
SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg487_out;
SharedReg861_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg861_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg485_out;
SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1116_out;
SharedReg869_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg869_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg485_out;
SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1116_out;
SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg855_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg484_out;
SharedReg294_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg294_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg484_out;
SharedReg486_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg486_out;
SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg295_out;
SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg295_out;
SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg860_out;
SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg860_out;
SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg677_out;
SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg489_out;
SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg488_out;
SharedReg1119_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1119_out;
SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg489_out;
SharedReg863_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg863_out;
SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg302_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg484_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg484_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg496_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg864_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1129_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg688_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg684_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1115_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg872_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1403_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg490_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1130_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg673_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg853_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1131_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg290_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg676_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg487_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg861_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg869_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg485_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1116_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg855_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg294_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg486_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg295_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg860_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg677_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1119_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg489_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg863_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg302_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg484_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg488_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No100_out);

SharedReg1119_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg676_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg676_out;
Delay37No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= Delay37No36_out;
SharedReg865_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg865_out;
Delay43No9_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= Delay43No9_out;
SharedReg496_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg496_out;
SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1117_out;
SharedReg1115_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1115_out;
SharedReg1127_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1127_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg673_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg484_out;
SharedReg1118_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1118_out;
SharedReg492_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg492_out;
SharedReg856_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg856_out;
SharedReg877_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg877_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg673_out;
SharedReg313_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg313_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg485_out;
SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg484_out;
SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg687_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg673_out;
SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1117_out;
SharedReg858_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg858_out;
SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg485_out;
SharedReg690_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg690_out;
SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg292_out;
SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg36_out;
SharedReg1404_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1404_out;
SharedReg499_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg499_out;
SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg290_out;
SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1120_out;
SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1120_out;
SharedReg881_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg881_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg673_out;
SharedReg1400_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1400_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg673_out;
SharedReg876_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg876_out;
SharedReg674_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg674_out;
SharedReg63_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg63_out;
SharedReg1116_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1116_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg673_out;
SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg290_out;
SharedReg854_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg854_out;
SharedReg1402_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1402_out;
SharedReg1126_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1126_out;
SharedReg1121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1121_out;
SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg675_out;
SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1117_out;
SharedReg689_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg689_out;
SharedReg853_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg853_out;
SharedReg37_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg37_out;
SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg675_out;
SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg675_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay37No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg865_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay43No9_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg496_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1115_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1127_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1118_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg492_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg856_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg877_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg313_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg484_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg687_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg858_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg485_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg690_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1404_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg499_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1120_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg881_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1400_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg876_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg674_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg63_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1116_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg290_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg854_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1402_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1126_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1117_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg689_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg853_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg37_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg675_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg676_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No102_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg509_out;
SharedReg1139_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1139_out;
SharedReg510_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg510_out;
SharedReg1410_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1410_out;
SharedReg77_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg505_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg8_out;
SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg509_out;
SharedReg517_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg517_out;
SharedReg893_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg893_out;
SharedReg1149_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1149_out;
SharedReg708_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg708_out;
SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg693_out;
SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg697_out;
SharedReg704_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg704_out;
SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg511_out;
SharedReg1136_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1136_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg505_out;
SharedReg1135_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1135_out;
SharedReg1418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1418_out;
SharedReg1350_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1350_out;
SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg506_out;
SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg322_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg505_out;
SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg511_out;
SharedReg1150_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1150_out;
SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg697_out;
SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg693_out;
SharedReg882_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg882_out;
SharedReg1151_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1151_out;
SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg506_out;
SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg317_out;
SharedReg329_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg329_out;
SharedReg884_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg884_out;
SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg508_out;
SharedReg82_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg82_out;
SharedReg696_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg696_out;
SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg508_out;
SharedReg890_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg890_out;
SharedReg897_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg897_out;
SharedReg76_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg76_out;
SharedReg83_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg83_out;
SharedReg883_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg883_out;
SharedReg319_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg319_out;
SharedReg68_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg68_out;
SharedReg701_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg701_out;
SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg527_out;
SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1156_out;
SharedReg926_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg926_out;
SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg527_out;
SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1156_out;
SharedReg1349_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1349_out;
SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg526_out;
SharedReg99_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg99_out;
SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg526_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1139_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg509_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg517_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg893_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1149_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg510_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg708_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg704_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1136_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1135_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1350_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1410_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg511_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1150_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg697_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg693_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg882_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1151_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg506_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg77_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg329_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg884_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg82_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg696_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg508_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg890_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg897_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg76_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg83_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg883_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg319_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg68_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg701_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg926_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg527_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1156_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1349_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg99_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg526_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg505_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No102_out);

SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg695_out;
SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg709_out;
SharedReg1400_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1400_out;
SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg695_out;
SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg695_out;
SharedReg1139_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1139_out;
SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
SharedReg696_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg696_out;
Delay37No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast <= Delay37No37_out;
SharedReg894_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg894_out;
Delay43No10_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast <= Delay43No10_out;
SharedReg517_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg517_out;
SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1135_out;
SharedReg1147_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1147_out;
SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg693_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg505_out;
SharedReg1138_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1138_out;
SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg513_out;
SharedReg885_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg885_out;
SharedReg905_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg905_out;
SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg693_out;
SharedReg339_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg339_out;
SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg506_out;
SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg505_out;
SharedReg707_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg707_out;
SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg693_out;
SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1137_out;
SharedReg887_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg887_out;
SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg506_out;
SharedReg710_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg710_out;
SharedReg319_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg319_out;
SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg66_out;
SharedReg1351_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1351_out;
SharedReg520_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg520_out;
SharedReg317_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg317_out;
SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1140_out;
SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1140_out;
SharedReg909_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg909_out;
SharedReg882_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg882_out;
SharedReg340_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg340_out;
SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg66_out;
SharedReg904_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg904_out;
SharedReg91_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg91_out;
SharedReg335_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg335_out;
SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1135_out;
SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg713_out;
SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg713_out;
SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg910_out;
SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg713_out;
SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg713_out;
SharedReg932_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg932_out;
SharedReg714_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg714_out;
SharedReg120_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg120_out;
SharedReg1156_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1156_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg696_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay37No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg894_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay43No10_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg709_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg517_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1147_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1138_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg513_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg885_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg905_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1400_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg339_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg505_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg707_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg693_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1137_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg887_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg710_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg319_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1351_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg520_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg317_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1140_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg909_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg882_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg340_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg66_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg904_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg91_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg335_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1135_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg713_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg695_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg932_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg714_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg120_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1156_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1139_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No104_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg956_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg956_out;
SharedReg548_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg548_out;
SharedReg1176_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1176_out;
SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg347_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg347_out;
SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg547_out;
SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg530_out;
SharedReg1159_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1159_out;
SharedReg531_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg531_out;
SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg892_out;
SharedReg329_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg329_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg526_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg526_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg526_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg8_out;
SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg530_out;
SharedReg538_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg538_out;
SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg921_out;
SharedReg1169_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1169_out;
SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg728_out;
SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg713_out;
SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg717_out;
SharedReg724_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg724_out;
SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg532_out;
SharedReg1156_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1156_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg526_out;
SharedReg1155_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1155_out;
SharedReg1364_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1364_out;
SharedReg1431_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1431_out;
SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg527_out;
SharedReg348_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg348_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg526_out;
SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg532_out;
SharedReg1170_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1170_out;
SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg717_out;
SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg713_out;
SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg910_out;
SharedReg1171_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1171_out;
SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg527_out;
SharedReg343_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg343_out;
SharedReg920_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg920_out;
SharedReg357_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg357_out;
SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg717_out;
SharedReg1437_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1437_out;
SharedReg721_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg721_out;
SharedReg352_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg352_out;
SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1436_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg380_out;
SharedReg1430_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1430_out;
SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg550_out;
SharedReg140_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg140_out;
SharedReg736_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg736_out;
SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg550_out;
SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1436_out;
SharedReg955_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg955_out;
SharedReg134_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg134_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg956_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg548_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg329_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1176_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg538_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1169_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg724_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1156_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1155_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1364_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1431_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg348_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg526_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg532_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1170_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg713_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1171_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg527_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg343_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg920_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg357_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg347_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg717_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1437_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg721_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg352_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1430_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg140_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg736_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg547_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg550_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1436_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg955_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg134_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg530_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1159_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg531_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No104_out);

SharedReg1428_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1428_out;
SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg733_out;
SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg733_out;
SharedReg962_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg962_out;
SharedReg734_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg734_out;
SharedReg149_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg149_out;
SharedReg1176_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1176_out;
SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg715_out;
SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1157_out;
SharedReg729_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg729_out;
SharedReg1347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1347_out;
SharedReg318_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg318_out;
SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg715_out;
SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg715_out;
SharedReg1159_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1159_out;
SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg26_out;
SharedReg716_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg716_out;
Delay37No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast <= Delay37No38_out;
SharedReg922_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg922_out;
Delay43No11_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast <= Delay43No11_out;
SharedReg538_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg538_out;
SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1157_out;
SharedReg1155_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1155_out;
SharedReg1167_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1167_out;
SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg713_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg526_out;
SharedReg1158_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1158_out;
SharedReg534_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg534_out;
SharedReg913_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg913_out;
SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg935_out;
SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg713_out;
SharedReg122_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg122_out;
SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg527_out;
SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg526_out;
SharedReg727_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg727_out;
SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg713_out;
SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1157_out;
SharedReg915_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg915_out;
SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg527_out;
SharedReg730_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg730_out;
SharedReg345_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg345_out;
SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg910_out;
SharedReg344_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg344_out;
SharedReg1173_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1173_out;
SharedReg919_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg919_out;
SharedReg728_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg728_out;
SharedReg123_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg123_out;
SharedReg936_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg936_out;
SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg343_out;
SharedReg1325_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1325_out;
SharedReg562_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg562_out;
SharedReg124_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg124_out;
SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1180_out;
SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1180_out;
SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg967_out;
SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg910_out;
SharedReg151_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg151_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1428_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg318_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1159_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg733_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg716_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay37No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg922_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay43No11_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg538_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1155_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg962_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1167_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1158_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg534_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg913_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg122_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg734_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg526_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg727_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg713_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg915_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg527_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg730_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg345_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg344_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg149_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1173_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg919_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg728_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg123_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg936_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1325_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg562_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg124_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1176_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1180_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg910_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg151_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg715_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1157_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg729_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No106_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg171_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg171_out;
SharedReg756_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg948_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg948_out;
SharedReg983_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg983_out;
SharedReg379_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg379_out;
SharedReg984_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg984_out;
SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg569_out;
SharedReg1196_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1196_out;
SharedReg942_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg942_out;
SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg568_out;
SharedReg372_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg372_out;
SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg568_out;
SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg551_out;
SharedReg1179_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1179_out;
SharedReg552_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg552_out;
SharedReg920_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg920_out;
SharedReg355_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg355_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg547_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg8_out;
SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg551_out;
SharedReg559_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg559_out;
SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg951_out;
SharedReg1189_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1189_out;
SharedReg748_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg748_out;
SharedReg733_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg733_out;
SharedReg737_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg737_out;
SharedReg744_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg744_out;
SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg553_out;
SharedReg1176_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1176_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg547_out;
SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1175_out;
SharedReg1445_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1445_out;
SharedReg1324_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1324_out;
SharedReg548_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg548_out;
SharedReg373_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg373_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg547_out;
SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg553_out;
SharedReg564_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg564_out;
SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1175_out;
SharedReg374_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg374_out;
SharedReg124_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg124_out;
SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg951_out;
SharedReg380_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg380_out;
SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg951_out;
SharedReg1210_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1210_out;
SharedReg757_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg757_out;
SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg753_out;
SharedReg1321_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1321_out;
SharedReg1211_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1211_out;
SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg569_out;
SharedReg368_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg368_out;
SharedReg978_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg978_out;
SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg410_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg942_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg372_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1179_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg552_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg920_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg355_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg756_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg571_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg551_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg559_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1189_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg748_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg733_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg737_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg744_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1176_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg948_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1445_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1324_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg548_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg373_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg547_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg553_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg564_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1175_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg983_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg374_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg124_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg380_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg951_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1210_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg757_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1321_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1211_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg379_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg368_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg978_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg984_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg569_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1196_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No106_out);

SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg583_out;
SharedReg368_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg368_out;
SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1200_out;
SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1200_out;
SharedReg997_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg997_out;
SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg940_out;
SharedReg393_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg393_out;
SharedReg1321_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1321_out;
SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg753_out;
SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg753_out;
SharedReg992_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg992_out;
SharedReg754_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg754_out;
SharedReg391_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg391_out;
SharedReg1196_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1196_out;
SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg735_out;
SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1177_out;
SharedReg749_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg749_out;
SharedReg1428_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1428_out;
SharedReg344_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg344_out;
SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg735_out;
SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg735_out;
SharedReg1179_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1179_out;
SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg26_out;
SharedReg736_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg736_out;
Delay37No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast <= Delay37No39_out;
SharedReg952_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg952_out;
Delay43No12_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast <= Delay43No12_out;
SharedReg559_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg559_out;
SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1177_out;
SharedReg1175_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1175_out;
SharedReg1187_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1187_out;
SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg733_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg547_out;
SharedReg1178_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1178_out;
SharedReg555_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg555_out;
SharedReg943_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg943_out;
SharedReg1453_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1453_out;
SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg733_out;
SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg364_out;
SharedReg548_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg548_out;
SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg547_out;
SharedReg1188_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1188_out;
SharedReg1181_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1181_out;
SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg369_out;
SharedReg374_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg374_out;
SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg940_out;
SharedReg124_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg124_out;
SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg940_out;
SharedReg767_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg767_out;
SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg753_out;
SharedReg1197_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1197_out;
SharedReg1326_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1326_out;
SharedReg569_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg569_out;
SharedReg770_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg770_out;
SharedReg156_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg156_out;
SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg940_out;
SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg369_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg368_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg992_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg754_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg391_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1196_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg749_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1428_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg344_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg735_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1179_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1200_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg736_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => Delay37No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg952_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay43No12_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg559_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1177_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1175_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1187_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg997_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1178_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg555_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg943_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1453_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg733_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg364_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg548_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg547_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1188_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1181_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg374_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg124_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg767_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1197_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1326_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg569_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg393_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg770_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg156_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg940_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg369_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1321_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg753_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No108_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg773_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg773_out;
SharedReg968_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg968_out;
SharedReg1231_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1231_out;
SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg590_out;
SharedReg154_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg1008_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1008_out;
SharedReg196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg196_out;
SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg592_out;
SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg412_out;
SharedReg776_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg592_out;
SharedReg1329_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1329_out;
SharedReg1015_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1015_out;
SharedReg165_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg165_out;
SharedReg1016_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1016_out;
SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg590_out;
SharedReg1216_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1216_out;
SharedReg970_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg970_out;
SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg589_out;
SharedReg400_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg400_out;
SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg589_out;
SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg572_out;
SharedReg1199_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1199_out;
SharedReg573_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg573_out;
SharedReg950_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg950_out;
SharedReg380_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg380_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg568_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg8_out;
SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg572_out;
SharedReg580_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg580_out;
SharedReg979_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg979_out;
SharedReg1209_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1209_out;
SharedReg768_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg768_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg753_out;
SharedReg757_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg757_out;
SharedReg764_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg764_out;
SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg574_out;
SharedReg1196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1196_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg568_out;
SharedReg386_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg386_out;
SharedReg959_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg959_out;
SharedReg158_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg158_out;
SharedReg1195_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1195_out;
SharedReg971_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg971_out;
SharedReg144_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg144_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg753_out;
SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1215_out;
SharedReg1018_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1018_out;
SharedReg1030_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1030_out;
SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg590_out;
SharedReg188_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg188_out;
SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg589_out;
SharedReg595_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg595_out;
SharedReg606_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg606_out;
SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1215_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg773_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg968_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1329_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1015_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg165_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1016_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1216_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg970_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg400_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1231_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1199_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg573_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg950_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg380_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg580_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg979_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg154_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1209_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg768_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg757_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg764_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg386_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg959_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1008_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg158_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1195_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg971_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg144_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1018_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1030_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg590_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg188_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg196_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg589_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg595_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg606_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1215_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg592_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No108_out);

SharedReg1217_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1217_out;
SharedReg973_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg973_out;
SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg590_out;
SharedReg790_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg790_out;
SharedReg398_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg398_out;
SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg397_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg397_out;
SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg604_out;
SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg396_out;
SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1220_out;
SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1220_out;
SharedReg1056_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1056_out;
SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg968_out;
SharedReg423_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg423_out;
SharedReg998_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg998_out;
SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg773_out;
SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg773_out;
SharedReg1051_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1051_out;
SharedReg774_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg774_out;
SharedReg421_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg421_out;
SharedReg1216_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1216_out;
SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg755_out;
SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1197_out;
SharedReg769_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg769_out;
SharedReg1321_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1321_out;
SharedReg369_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg369_out;
SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg755_out;
SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg755_out;
SharedReg1199_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1199_out;
SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg26_out;
SharedReg756_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg756_out;
Delay37No40_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast <= Delay37No40_out;
SharedReg980_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg980_out;
Delay43No13_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast <= Delay43No13_out;
SharedReg580_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg580_out;
SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1197_out;
SharedReg1195_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1195_out;
SharedReg1207_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1207_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg753_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg568_out;
SharedReg1198_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1198_out;
SharedReg370_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg370_out;
SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1001_out;
SharedReg150_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg150_out;
SharedReg1206_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1206_out;
SharedReg1345_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1345_out;
SharedReg162_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg162_out;
SharedReg1200_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1200_out;
SharedReg597_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg597_out;
SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1001_out;
SharedReg993_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg993_out;
SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg773_out;
SharedReg422_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg422_out;
SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg590_out;
SharedReg589_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg589_out;
SharedReg1228_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1228_out;
SharedReg1221_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1221_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1217_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg973_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1056_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg423_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg998_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1051_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg774_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg421_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1216_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg769_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1321_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg369_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg755_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1199_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg790_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg756_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => Delay37No40_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg980_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg398_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => Delay43No13_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg580_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1197_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1195_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1207_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg568_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1198_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg370_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg968_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg150_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1206_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1345_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg162_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1200_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg597_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1001_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg993_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg773_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg422_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg397_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg590_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg589_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1228_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1221_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1220_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Subtract2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_5_impl_out,
                 X => Delay1No110_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg189_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg154_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1009_out;
SharedReg194_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1009_out;
SharedReg1250_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1250_out;
SharedReg797_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg797_out;
SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg777_out;
SharedReg1007_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1007_out;
SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg781_out;
SharedReg405_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg976_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg976_out;
SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg438_out;
SharedReg1000_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1000_out;
SharedReg413_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg413_out;
SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg969_out;
SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg398_out;
SharedReg156_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg156_out;
SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg781_out;
SharedReg611_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg611_out;
SharedReg1236_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1236_out;
SharedReg591_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg591_out;
SharedReg401_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg401_out;
SharedReg159_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg159_out;
SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1328_out;
SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1328_out;
SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg777_out;
SharedReg594_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg594_out;
SharedReg1195_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1195_out;
SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg13_out;
SharedReg385_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg385_out;
SharedReg957_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg957_out;
SharedReg165_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg165_out;
SharedReg766_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg766_out;
SharedReg1208_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1208_out;
SharedReg577_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg577_out;
SharedReg396_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg396_out;
SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg969_out;
SharedReg968_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg968_out;
SharedReg999_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg999_out;
SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg398_out;
SharedReg788_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg788_out;
SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg773_out;
SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg777_out;
SharedReg784_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg784_out;
SharedReg595_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg595_out;
SharedReg1216_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1216_out;
SharedReg589_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg589_out;
SharedReg415_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg415_out;
SharedReg987_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg987_out;
SharedReg187_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg187_out;
SharedReg1215_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1215_out;
SharedReg1001_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1001_out;
SharedReg175_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg175_out;
SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg773_out;
SharedReg1235_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1235_out;
SharedReg1392_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1392_out;
   MUX_Subtract2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg976_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1000_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg413_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg156_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg611_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1236_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg591_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg401_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg159_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1328_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg594_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1195_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg194_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg17_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg13_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg385_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg957_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg165_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1009_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg766_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1208_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg577_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg396_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg969_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg968_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg999_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg398_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg788_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1250_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg784_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg595_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1216_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg589_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg415_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg987_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg187_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1215_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1001_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg797_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg175_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg773_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1235_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1392_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg777_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1007_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg781_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_5_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_0_out,
                 Y => Delay1No110_out);

SharedReg397_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg189_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg968_out;
SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg154_out;
SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg968_out;
SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg807_out;
SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg793_out;
SharedReg1233_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1233_out;
SharedReg977_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg977_out;
SharedReg788_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg788_out;
SharedReg209_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg209_out;
SharedReg994_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg994_out;
SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg183_out;
SharedReg1377_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1377_out;
SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg154_out;
SharedReg1051_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1051_out;
SharedReg207_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg207_out;
SharedReg445_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg445_out;
SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1215_out;
SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg793_out;
SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg793_out;
SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg773_out;
SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg396_out;
SharedReg969_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg969_out;
SharedReg1000_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1000_out;
SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1226_out;
SharedReg1221_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1221_out;
SharedReg1198_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1198_out;
SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg31_out;
SharedReg380_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg380_out;
SharedReg1334_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1334_out;
SharedReg167_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg167_out;
Delay41No22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast <= Delay41No22_out;
SharedReg1211_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1211_out;
SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg765_out;
SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg169_out;
SharedReg982_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg982_out;
SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg996_out;
SharedReg1026_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1026_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg425_out;
SharedReg601_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg601_out;
SharedReg1217_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1217_out;
SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1215_out;
SharedReg1227_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1227_out;
SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg773_out;
SharedReg589_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg589_out;
SharedReg1218_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1218_out;
SharedReg398_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg398_out;
SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1030_out;
SharedReg181_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg181_out;
SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1226_out;
SharedReg1025_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1025_out;
SharedReg191_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg191_out;
SharedReg1220_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1220_out;
SharedReg618_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg618_out;
SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1030_out;
   MUX_Subtract2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg209_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg994_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1377_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1051_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg207_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg445_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg396_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg969_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1000_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1221_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1198_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg154_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg35_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg31_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg380_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1334_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg167_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg968_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => Delay41No22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1211_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg982_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1026_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg601_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1217_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1215_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1227_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg773_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg589_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1218_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg398_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg181_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1226_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1025_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg793_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg191_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1220_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg618_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1030_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1233_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg977_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg788_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_5_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Subtract2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_6_impl_out,
                 X => Delay1No112_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1376_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1376_out;
SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg611_out;
SharedReg431_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg431_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg610_out;
SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg616_out;
SharedReg627_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg627_out;
SharedReg1235_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1235_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg793_out;
SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1027_out;
SharedReg1251_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1251_out;
SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg611_out;
SharedReg183_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg183_out;
SharedReg1036_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1036_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg440_out;
SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg613_out;
SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg200_out;
SharedReg796_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg796_out;
SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg613_out;
SharedReg1006_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1006_out;
SharedReg1042_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1042_out;
SharedReg193_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg193_out;
SharedReg1043_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1043_out;
SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg611_out;
SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1236_out;
SharedReg1029_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1029_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg610_out;
SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg430_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg610_out;
SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg593_out;
SharedReg1219_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1219_out;
SharedReg594_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg594_out;
SharedReg978_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg978_out;
SharedReg408_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg408_out;
SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg589_out;
SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg589_out;
SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg589_out;
SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg8_out;
SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg593_out;
SharedReg601_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg601_out;
SharedReg1037_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1037_out;
SharedReg1229_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1229_out;
SharedReg1228_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1228_out;
SharedReg598_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg598_out;
SharedReg426_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg426_out;
SharedReg1028_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1028_out;
SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1027_out;
SharedReg1374_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1374_out;
SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg428_out;
SharedReg808_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg808_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg793_out;
SharedReg797_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg797_out;
SharedReg804_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg804_out;
SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg616_out;
SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1236_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg610_out;
SharedReg444_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg444_out;
SharedReg1046_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1046_out;
   MUX_Subtract2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1376_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg183_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1036_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg796_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg613_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1006_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1042_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg431_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg193_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1043_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg611_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1029_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1219_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg594_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg978_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg408_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg589_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg14_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg593_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg601_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1037_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1229_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1228_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg598_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg627_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg426_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1028_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1374_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg808_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg797_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg804_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg616_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1235_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1236_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg610_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg444_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1046_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg793_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1027_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1251_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_6_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_0_out,
                 Y => Delay1No112_out);

SharedReg1052_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1052_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg793_out;
SharedReg451_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg611_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg610_out;
SharedReg1248_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1248_out;
SharedReg1241_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1241_out;
SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1237_out;
SharedReg1003_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1003_out;
SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg611_out;
SharedReg810_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg810_out;
SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg428_out;
SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1027_out;
SharedReg427_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg427_out;
SharedReg625_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg625_out;
SharedReg426_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg426_out;
SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1240_out;
SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1240_out;
SharedReg1399_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1399_out;
SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1027_out;
SharedReg452_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg452_out;
SharedReg1373_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1373_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg793_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg793_out;
SharedReg1080_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1080_out;
SharedReg794_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg794_out;
SharedReg450_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg450_out;
SharedReg1236_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1236_out;
SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg775_out;
SharedReg1217_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1217_out;
SharedReg789_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg789_out;
SharedReg998_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg998_out;
SharedReg397_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg397_out;
SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg775_out;
SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg775_out;
SharedReg1219_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1219_out;
SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg26_out;
SharedReg776_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg776_out;
Delay37No41_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast <= Delay37No41_out;
SharedReg1039_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1039_out;
Delay43No14_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast <= Delay43No14_out;
SharedReg1231_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1231_out;
SharedReg785_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg785_out;
SharedReg198_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg198_out;
SharedReg1041_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1041_out;
SharedReg1055_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1055_out;
SharedReg1398_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1398_out;
SharedReg454_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg454_out;
SharedReg622_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg622_out;
SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1237_out;
SharedReg1235_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1235_out;
SharedReg1247_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1247_out;
SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg793_out;
SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg610_out;
SharedReg1238_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1238_out;
SharedReg185_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg185_out;
SharedReg1376_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1376_out;
   MUX_Subtract2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1052_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg810_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg427_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg625_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg426_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1240_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1399_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1027_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg451_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg452_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1373_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1080_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg794_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg450_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1236_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1217_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg789_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg998_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg397_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg775_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1219_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg32_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg25_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg776_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => Delay37No41_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1039_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => Delay43No14_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1231_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg785_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1248_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg198_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1041_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1055_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1398_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg454_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg622_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1235_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1247_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg793_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1241_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg610_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1238_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg185_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1376_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1237_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1003_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg611_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_6_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Subtract2_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_7_impl_out,
                 X => Delay1No114_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast);

SharedReg817_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg817_out;
SharedReg824_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg824_out;
SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg637_out;
SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1256_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg631_out;
SharedReg253_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg253_out;
SharedReg1076_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1076_out;
SharedReg1060_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1060_out;
SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg632_out;
SharedReg215_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg215_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg631_out;
SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg637_out;
SharedReg648_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg648_out;
SharedReg1255_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1255_out;
SharedReg813_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg813_out;
SharedReg1057_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1057_out;
SharedReg1271_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1271_out;
SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg632_out;
SharedReg210_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg210_out;
SharedReg1066_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1066_out;
SharedReg249_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg249_out;
SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg634_out;
SharedReg442_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg442_out;
SharedReg816_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg816_out;
SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg634_out;
SharedReg1381_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1381_out;
SharedReg1074_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1074_out;
SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg220_out;
SharedReg1390_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1390_out;
SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg632_out;
SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1256_out;
SharedReg1059_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1059_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg631_out;
SharedReg239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg239_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg631_out;
SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg614_out;
SharedReg1239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1239_out;
SharedReg615_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg615_out;
SharedReg1036_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1036_out;
SharedReg438_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg438_out;
SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg610_out;
SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg610_out;
SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg610_out;
SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg13_out;
SharedReg443_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg443_out;
SharedReg1044_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1044_out;
SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg220_out;
SharedReg806_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg806_out;
SharedReg10_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg8_out;
SharedReg635_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg635_out;
SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg643_out;
SharedReg1097_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1097_out;
SharedReg1269_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1269_out;
SharedReg1268_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1268_out;
SharedReg640_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg640_out;
   MUX_Subtract2_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg817_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg824_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg648_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1255_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg813_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1057_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1271_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg210_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1066_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg637_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg249_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg442_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg816_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg634_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1381_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1074_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1390_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1256_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1059_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1239_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg615_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1036_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg438_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg631_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg610_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg2_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg14_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg12_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg16_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg253_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg13_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg443_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1044_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg220_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg806_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg10_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg9_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg8_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg635_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1076_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1097_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1269_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1268_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg640_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1060_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg632_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg215_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_7_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_7_impl_0_out,
                 Y => Delay1No114_out);

SharedReg1255_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1255_out;
SharedReg1267_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1267_out;
SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg813_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg631_out;
SharedReg1258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1258_out;
SharedReg428_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg428_out;
SharedReg1060_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1060_out;
SharedReg1081_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1081_out;
SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg813_out;
SharedReg257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg257_out;
SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg632_out;
SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg631_out;
SharedReg1268_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1268_out;
SharedReg1261_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1261_out;
SharedReg1257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1257_out;
SharedReg1378_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1378_out;
SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg632_out;
SharedReg830_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg830_out;
SharedReg237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg237_out;
SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1057_out;
SharedReg236_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg236_out;
SharedReg646_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg646_out;
SharedReg235_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg235_out;
SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1260_out;
SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1260_out;
SharedReg1085_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1085_out;
SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1057_out;
SharedReg258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg258_out;
SharedReg1295_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1295_out;
SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg813_out;
SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg813_out;
SharedReg1317_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1317_out;
SharedReg814_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg814_out;
SharedReg256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg256_out;
SharedReg1256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1256_out;
SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg795_out;
SharedReg1237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1237_out;
SharedReg809_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg809_out;
SharedReg1373_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1373_out;
SharedReg427_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg427_out;
SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg795_out;
SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg795_out;
SharedReg1239_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1239_out;
SharedReg18_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_48_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg31_out;
SharedReg194_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg194_out;
SharedReg1386_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1386_out;
SharedReg222_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg222_out;
Delay41No24_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_55_cast <= Delay41No24_out;
SharedReg28_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg26_out;
SharedReg816_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg816_out;
Delay37No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_60_cast <= Delay37No43_out;
SharedReg1099_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1099_out;
Delay43No16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_62_cast <= Delay43No16_out;
SharedReg1271_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1271_out;
SharedReg825_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg825_out;
   MUX_Subtract2_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1255_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1267_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1268_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1261_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1378_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg632_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg830_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg236_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg646_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg235_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1260_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1085_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1057_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1295_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg631_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1317_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg814_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1256_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1237_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg809_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1373_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg427_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1258_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg795_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1239_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg18_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg32_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg25_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg30_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg428_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg31_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg194_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1386_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg222_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay41No24_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg28_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg27_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg26_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg816_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => Delay37No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1060_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1099_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => Delay43No16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1271_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg825_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1081_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg813_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg257_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_7_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_7_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Subtract2_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_8_impl_out,
                 X => Delay1No116_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg656_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg656_out;
SharedReg664_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg664_out;
SharedReg1466_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1466_out;
SharedReg846_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg846_out;
SharedReg1288_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1288_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg833_out;
SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg844_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg844_out;
SharedReg658_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg658_out;
SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1276_out;
SharedReg263_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg263_out;
SharedReg474_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg474_out;
SharedReg1473_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1473_out;
SharedReg1460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1460_out;
SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg653_out;
SharedReg461_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg461_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg652_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg833_out;
SharedReg669_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg669_out;
SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg837_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg833_out;
SharedReg1086_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1086_out;
SharedReg1291_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1291_out;
SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg653_out;
SharedReg1097_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1097_out;
SharedReg1305_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1305_out;
SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1088_out;
SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg655_out;
SharedReg279_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg279_out;
SharedReg836_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg836_out;
SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg655_out;
SharedReg1094_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1094_out;
SharedReg1102_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1102_out;
SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1276_out;
SharedReg1103_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1103_out;
SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg653_out;
SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1276_out;
SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1088_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg652_out;
SharedReg460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg460_out;
SharedReg635_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg635_out;
SharedReg1259_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1259_out;
SharedReg636_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg636_out;
SharedReg1066_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1066_out;
SharedReg247_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg247_out;
SharedReg631_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg631_out;
SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg837_out;
SharedReg1255_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1255_out;
SharedReg1_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg11_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg652_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg652_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg652_out;
SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_62_cast <= SharedReg4_out;
SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_63_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_64_cast <= SharedReg12_out;
   MUX_Subtract2_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg658_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg263_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg474_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1473_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg461_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg656_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg669_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1086_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1291_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1097_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1305_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg664_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg279_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg836_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg655_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1094_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1102_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1103_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg653_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1276_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1088_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1466_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg460_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg635_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1259_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg636_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1066_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg247_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg631_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1255_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg846_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg3_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg17_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg652_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg2_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1288_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg14_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg11_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg12_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg833_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg844_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_8_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_8_impl_0_out,
                 Y => Delay1No116_out);

SharedReg27_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg836_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg836_out;
Delay37No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast <= Delay37No44_out;
SharedReg1468_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1468_out;
Delay41No26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast <= Delay41No26_out;
SharedReg1291_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1291_out;
SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1277_out;
SharedReg1275_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1275_out;
SharedReg1287_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1287_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg833_out;
SharedReg652_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg652_out;
SharedReg483_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg483_out;
SharedReg237_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg237_out;
SharedReg1298_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1298_out;
SharedReg1110_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1110_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg833_out;
SharedReg480_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg480_out;
SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg653_out;
SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1280_out;
SharedReg1288_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1288_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg833_out;
SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1277_out;
SharedReg1300_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1300_out;
SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg653_out;
SharedReg850_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg850_out;
SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1457_out;
SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1086_out;
SharedReg1090_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1090_out;
SharedReg667_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg667_out;
SharedReg457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg457_out;
SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1280_out;
SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1280_out;
SharedReg1111_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1111_out;
SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1086_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg833_out;
SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1457_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg833_out;
SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg833_out;
SharedReg1109_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1109_out;
SharedReg834_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg834_out;
SharedReg285_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg285_out;
SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg815_out;
SharedReg1257_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1257_out;
SharedReg829_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg829_out;
SharedReg1295_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1295_out;
SharedReg236_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg236_out;
SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg815_out;
SharedReg1286_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1286_out;
SharedReg1258_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1258_out;
SharedReg19_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_55_cast <= SharedReg29_out;
SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg835_out;
SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg835_out;
SharedReg1279_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1279_out;
SharedReg18_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_62_cast <= SharedReg22_out;
SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_63_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_64_cast <= SharedReg30_out;
   MUX_Subtract2_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg652_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg483_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg237_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1298_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1110_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg480_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg836_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1288_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1300_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg653_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg850_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1090_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg667_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => Delay37No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1280_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1111_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1086_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1457_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg833_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1109_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1468_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg834_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg285_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1257_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg829_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1295_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg236_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg815_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1286_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1258_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => Delay41No26_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg19_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg21_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg35_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg24_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg835_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1279_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg18_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1291_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg32_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg29_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg30_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1277_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1275_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1287_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_8_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_8_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No118_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1584_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1612_out;
SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg854_out;
SharedReg1536_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1536_out;
SharedReg1423_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1423_out;
SharedReg1400_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1400_out;
SharedReg1650_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1650_out;
SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg1484_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1539_out;
SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1404_out;
SharedReg295_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg295_out;
SharedReg1589_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1647_out;
SharedReg299_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg299_out;
SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg43_out;
SharedReg1491_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1493_out;
SharedReg302_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg302_out;
SharedReg1495_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1629_out;
SharedReg303_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg303_out;
SharedReg1414_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1414_out;
SharedReg1577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1577_out;
SharedReg1412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1412_out;
SharedReg1529_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1590_out;
SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg853_out;
SharedReg1598_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1505_out;
SharedReg1408_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1408_out;
SharedReg858_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg858_out;
SharedReg1558_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1558_out;
SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg44_out;
SharedReg1645_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1645_out;
SharedReg859_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg859_out;
SharedReg1619_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1607_out;
SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1404_out;
SharedReg1530_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1608_out;
SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg853_out;
SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg853_out;
SharedReg1609_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1611_out;
SharedReg1421_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1421_out;
SharedReg1534_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1534_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1584_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1626_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1539_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg295_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1589_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1488_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1649_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1647_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg299_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1491_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1612_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1545_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1602_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1493_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg302_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1495_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1548_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1549_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1614_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1629_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg303_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg854_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1414_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1412_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1529_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1579_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1642_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1596_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1590_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1598_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1536_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1592_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1637_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1505_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1408_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg858_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1558_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1645_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg859_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1619_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1423_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1606_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1607_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1404_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1530_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1580_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1608_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg853_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1609_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1624_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1400_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1610_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1611_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1421_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1534_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1650_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1484_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No118_out);

SharedReg874_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg874_out;
SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg853_out;
SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg854_out;
SharedReg1627_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1627_out;
SharedReg1422_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1422_out;
SharedReg1587_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1537_out;
SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1400_out;
SharedReg1538_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1538_out;
SharedReg290_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg290_out;
SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg1651_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1540_out;
SharedReg857_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg857_out;
SharedReg1408_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1408_out;
SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1403_out;
SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1404_out;
SharedReg1543_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1544_out;
SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg865_out;
SharedReg45_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg45_out;
SharedReg864_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg864_out;
SharedReg304_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg304_out;
SharedReg1546_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1546_out;
SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg47_out;
SharedReg305_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg305_out;
SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg48_out;
SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1413_out;
SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1413_out;
SharedReg1575_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1576_out;
SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg49_out;
SharedReg1578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1578_out;
SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1413_out;
SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg48_out;
SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg853_out;
SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1400_out;
SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1401_out;
SharedReg1643_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1643_out;
SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1400_out;
SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1401_out;
SharedReg856_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg856_out;
SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg40_out;
SharedReg1644_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1557_out;
SharedReg1407_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1407_out;
SharedReg1559_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1559_out;
SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg860_out;
SharedReg1618_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1618_out;
SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1403_out;
SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1404_out;
SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1403_out;
SharedReg1620_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1620_out;
SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg55_out;
SharedReg1420_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1420_out;
SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg860_out;
SharedReg1622_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1623_out;
SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg854_out;
SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg853_out;
SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg854_out;
SharedReg858_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg858_out;
SharedReg1582_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1582_out;
SharedReg312_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg312_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg874_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1651_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1540_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg857_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1408_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1543_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1544_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg865_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg45_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg864_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg304_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1546_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg305_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1575_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1627_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1576_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1413_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1643_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1422_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1401_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg856_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1644_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1557_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1407_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1559_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1618_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1587_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1404_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1403_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1620_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg55_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1420_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg860_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1622_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1623_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg853_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1537_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg854_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg858_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1582_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg312_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1400_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1538_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg290_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No120_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1400_out;
SharedReg1609_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1611_out;
SharedReg1366_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1366_out;
SharedReg1534_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1612_out;
SharedReg883_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg883_out;
SharedReg1536_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1536_out;
SharedReg1368_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1368_out;
SharedReg1347_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1347_out;
SharedReg1650_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1650_out;
SharedReg66_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg66_out;
SharedReg1484_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1539_out;
SharedReg1351_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1351_out;
SharedReg322_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg322_out;
SharedReg1589_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1647_out;
SharedReg326_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg326_out;
SharedReg73_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg73_out;
SharedReg1491_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1493_out;
SharedReg329_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg329_out;
SharedReg1495_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1629_out;
SharedReg330_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg330_out;
SharedReg1361_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1361_out;
SharedReg1577_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1577_out;
SharedReg1359_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1359_out;
SharedReg1529_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1590_out;
SharedReg882_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg882_out;
SharedReg1598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1505_out;
SharedReg1355_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1355_out;
SharedReg887_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg887_out;
SharedReg1558_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1558_out;
SharedReg74_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg74_out;
SharedReg1645_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1645_out;
SharedReg888_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg888_out;
SharedReg1619_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1607_out;
SharedReg886_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg886_out;
SharedReg1530_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1608_out;
SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1400_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1609_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg883_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1536_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1368_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1347_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1650_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg66_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1484_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1539_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1351_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg322_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1624_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1589_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1488_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1649_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1647_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg326_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg73_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1491_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1545_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1602_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1493_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1610_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg329_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1495_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1548_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1549_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1614_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1629_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg330_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1361_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1577_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1359_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1611_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1529_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1579_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1642_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1596_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1590_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg882_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1592_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1637_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1505_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1366_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1355_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg887_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1558_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg74_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1645_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg888_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1619_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1606_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1607_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg886_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1534_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1530_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1580_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1608_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1400_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1584_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1626_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1612_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No120_out);

SharedReg1623_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1623_out;
SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1401_out;
SharedReg1400_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1400_out;
SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1401_out;
SharedReg1405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1405_out;
SharedReg1582_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1582_out;
SharedReg337_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg337_out;
SharedReg902_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg902_out;
SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg882_out;
SharedReg883_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg883_out;
SharedReg1627_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1627_out;
SharedReg1367_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1367_out;
SharedReg1587_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1537_out;
SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1347_out;
SharedReg1538_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1538_out;
SharedReg317_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg317_out;
SharedReg67_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg67_out;
SharedReg1651_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1540_out;
SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg886_out;
SharedReg1355_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1355_out;
SharedReg1350_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1350_out;
SharedReg1351_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1351_out;
SharedReg1543_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1544_out;
SharedReg894_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg894_out;
SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg75_out;
SharedReg893_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg893_out;
SharedReg331_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg331_out;
SharedReg1546_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1546_out;
SharedReg77_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg77_out;
SharedReg332_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg332_out;
SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg78_out;
SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1360_out;
SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1360_out;
SharedReg1575_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1576_out;
SharedReg79_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg79_out;
SharedReg1578_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1578_out;
SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1360_out;
SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg78_out;
SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg882_out;
SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1347_out;
SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1348_out;
SharedReg1643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1643_out;
SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1347_out;
SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1348_out;
SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg885_out;
SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg70_out;
SharedReg1644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1557_out;
SharedReg1354_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1354_out;
SharedReg1559_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1559_out;
SharedReg889_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg889_out;
SharedReg1618_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1618_out;
SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg886_out;
SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg885_out;
SharedReg1620_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1620_out;
SharedReg85_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg85_out;
SharedReg1365_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1365_out;
SharedReg1407_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1407_out;
SharedReg1622_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1622_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1623_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1627_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1367_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1587_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1537_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1538_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg317_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg67_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1651_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1540_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1400_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1355_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1350_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1351_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1543_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1544_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg894_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg893_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg331_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1401_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1546_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg77_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg332_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1575_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1576_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg79_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1578_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1405_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1360_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg78_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1347_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1348_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1582_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1557_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1354_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1559_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg889_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1618_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg886_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg885_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1620_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg337_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg85_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1365_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1407_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1622_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg902_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg882_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg883_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No122_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1606_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1607_out;
SharedReg1351_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1351_out;
SharedReg1530_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1608_out;
SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1347_out;
SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1347_out;
SharedReg1609_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1611_out;
SharedReg1447_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1447_out;
SharedReg1534_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1612_out;
SharedReg911_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg911_out;
SharedReg1536_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1536_out;
SharedReg1449_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1449_out;
SharedReg1428_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1428_out;
SharedReg1650_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1650_out;
SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg95_out;
SharedReg1484_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1539_out;
SharedReg1432_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1432_out;
SharedReg348_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg348_out;
SharedReg1589_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1647_out;
SharedReg352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg352_out;
SharedReg102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg102_out;
SharedReg1491_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1493_out;
SharedReg355_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg355_out;
SharedReg1495_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1629_out;
SharedReg356_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg356_out;
SharedReg1442_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1442_out;
SharedReg1577_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1577_out;
SharedReg1440_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1440_out;
SharedReg1529_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1590_out;
SharedReg910_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg910_out;
SharedReg1598_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1505_out;
SharedReg1436_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1436_out;
SharedReg1352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1352_out;
SharedReg1558_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1558_out;
SharedReg103_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg103_out;
SharedReg1645_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1645_out;
SharedReg1353_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1353_out;
SharedReg1619_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1619_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1606_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1607_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1610_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1611_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1447_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1534_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1584_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1626_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1612_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg911_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1536_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1449_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1351_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1428_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1650_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1484_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1539_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1432_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg348_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1589_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1488_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1649_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1530_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1647_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1491_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1545_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1602_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1493_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg355_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1495_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1548_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1580_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1549_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1614_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1629_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg356_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1442_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1577_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1440_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1529_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1579_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1642_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1608_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1596_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1590_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg910_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1598_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1592_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1637_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1505_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1436_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1352_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1558_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg103_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1645_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1353_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1619_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1347_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1609_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1624_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No122_out);

SharedReg1351_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1351_out;
SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1350_out;
SharedReg1620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1620_out;
SharedReg113_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg113_out;
SharedReg1446_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1446_out;
SharedReg889_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg889_out;
SharedReg1622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1623_out;
SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1348_out;
SharedReg1347_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1347_out;
SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1348_out;
SharedReg1352_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1352_out;
SharedReg1582_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1582_out;
SharedReg363_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg363_out;
SharedReg930_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg930_out;
SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg910_out;
SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg911_out;
SharedReg1627_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1627_out;
SharedReg1448_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1448_out;
SharedReg1587_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1537_out;
SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1428_out;
SharedReg1538_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1538_out;
SharedReg343_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg343_out;
SharedReg96_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg96_out;
SharedReg1651_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1540_out;
SharedReg914_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg914_out;
SharedReg1436_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1436_out;
SharedReg1431_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1431_out;
SharedReg1432_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1432_out;
SharedReg1543_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1544_out;
SharedReg922_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg922_out;
SharedReg104_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg104_out;
SharedReg921_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg921_out;
SharedReg357_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg357_out;
SharedReg1546_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1546_out;
SharedReg106_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg106_out;
SharedReg358_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg358_out;
SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg107_out;
SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1441_out;
SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1441_out;
SharedReg1575_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1576_out;
SharedReg108_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg108_out;
SharedReg1578_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1578_out;
SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1441_out;
SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg107_out;
SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg910_out;
SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1428_out;
SharedReg1429_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1429_out;
SharedReg1643_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1643_out;
SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg910_out;
SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg911_out;
SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg913_out;
SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg99_out;
SharedReg1644_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1557_out;
SharedReg1435_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1435_out;
SharedReg1559_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1559_out;
SharedReg1354_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1354_out;
SharedReg1618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1618_out;
SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1350_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1351_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1352_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1582_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg363_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg930_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1627_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1448_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1587_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1537_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1538_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg343_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg96_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1651_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg914_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1436_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1431_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg113_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1432_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1543_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1544_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg922_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg104_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg921_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg357_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1546_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg106_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg358_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1446_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1575_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg108_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1578_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1441_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg107_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg889_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1428_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1429_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1643_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg910_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1644_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1557_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1435_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1559_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1354_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1350_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1623_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1348_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1347_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No124_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg948_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg948_out;
SharedReg915_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg915_out;
SharedReg1558_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1558_out;
SharedReg351_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg351_out;
SharedReg1645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1645_out;
SharedReg916_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
SharedReg1619_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1607_out;
SharedReg1432_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1432_out;
SharedReg1530_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1608_out;
SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1428_out;
SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1428_out;
SharedReg1609_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1611_out;
SharedReg1340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1340_out;
SharedReg1534_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1612_out;
SharedReg941_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg941_out;
SharedReg1536_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1536_out;
SharedReg1342_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1342_out;
SharedReg1321_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1321_out;
SharedReg1650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1650_out;
SharedReg124_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg124_out;
SharedReg1484_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1539_out;
SharedReg1325_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1325_out;
SharedReg373_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg373_out;
SharedReg1589_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1647_out;
SharedReg377_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg377_out;
SharedReg350_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg350_out;
SharedReg1491_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1493_out;
SharedReg135_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg135_out;
SharedReg1495_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1629_out;
SharedReg381_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg381_out;
SharedReg1335_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1335_out;
SharedReg1577_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1577_out;
SharedReg1333_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1333_out;
SharedReg1529_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1590_out;
SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1428_out;
SharedReg1598_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1505_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg948_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg915_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1530_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1580_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1608_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1609_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1610_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1611_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1558_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1534_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1584_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1626_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1612_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg941_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1536_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1342_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1321_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg124_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg351_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1484_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1539_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1325_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg373_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1589_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1488_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1649_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1647_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg377_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg350_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1491_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1545_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1602_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1493_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg135_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1495_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1548_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1549_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1614_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1629_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg381_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1335_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1577_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1333_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1529_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1579_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1642_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1596_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1428_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1619_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1598_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1592_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1637_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1505_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1606_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1607_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1432_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No124_out);

SharedReg1644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1557_out;
SharedReg947_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg947_out;
SharedReg1559_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1559_out;
SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg1618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1618_out;
SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg913_out;
SharedReg914_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg914_out;
SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1431_out;
SharedReg1620_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1620_out;
SharedReg142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg142_out;
SharedReg1339_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1339_out;
SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg917_out;
SharedReg1622_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1623_out;
SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1429_out;
SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1428_out;
SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1429_out;
SharedReg1433_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1433_out;
SharedReg1582_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1582_out;
SharedReg389_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg389_out;
SharedReg960_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg960_out;
SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg941_out;
SharedReg1627_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1627_out;
SharedReg1341_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1341_out;
SharedReg1587_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1537_out;
SharedReg1321_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1321_out;
SharedReg1538_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1538_out;
SharedReg368_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg368_out;
SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg125_out;
SharedReg1651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1540_out;
SharedReg944_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg944_out;
SharedReg1329_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1329_out;
SharedReg1324_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1324_out;
SharedReg1325_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1325_out;
SharedReg1543_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1544_out;
SharedReg952_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg952_out;
SharedReg133_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg133_out;
SharedReg951_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg951_out;
SharedReg382_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg382_out;
SharedReg1546_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1546_out;
SharedReg135_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg135_out;
SharedReg383_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg383_out;
SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg136_out;
SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1334_out;
SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1334_out;
SharedReg1575_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1576_out;
SharedReg137_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg137_out;
SharedReg1578_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1578_out;
SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1334_out;
SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg136_out;
SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1428_out;
SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg941_out;
SharedReg1643_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1643_out;
SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1428_out;
SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1429_out;
SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1431_out;
SharedReg347_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg347_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1557_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1339_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1622_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1623_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1433_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1582_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg947_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg389_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg960_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1627_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1341_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1587_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1537_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1321_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1538_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1559_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg368_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1540_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg944_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1329_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1324_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1325_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1543_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1544_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg917_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg952_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg133_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg951_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg382_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1546_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg135_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg383_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1575_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1576_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg137_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1578_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1334_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg941_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1643_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1428_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1429_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg347_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg914_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1431_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1620_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No126_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1590_out;
SharedReg940_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg940_out;
SharedReg1598_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1505_out;
SharedReg1329_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1329_out;
SharedReg1433_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1433_out;
SharedReg1558_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1558_out;
SharedReg132_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg132_out;
SharedReg1645_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1645_out;
SharedReg946_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg946_out;
SharedReg1619_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1607_out;
SharedReg1325_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1325_out;
SharedReg1530_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1608_out;
SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1321_out;
SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1321_out;
SharedReg1609_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1611_out;
SharedReg988_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg988_out;
SharedReg1534_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1612_out;
SharedReg969_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg969_out;
SharedReg1536_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1536_out;
SharedReg990_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg990_out;
SharedReg998_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg998_out;
SharedReg1650_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1650_out;
SharedReg154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg154_out;
SharedReg1484_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1539_out;
SharedReg1002_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1002_out;
SharedReg401_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg401_out;
SharedReg1589_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1647_out;
SharedReg405_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg405_out;
SharedReg375_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg375_out;
SharedReg1491_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1493_out;
SharedReg166_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg166_out;
SharedReg1495_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1629_out;
SharedReg409_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg409_out;
SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1012_out;
SharedReg1577_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1577_out;
SharedReg1010_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1010_out;
SharedReg1529_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1642_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1590_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg132_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1645_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg946_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1619_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1606_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1607_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1325_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1530_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1580_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1608_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg940_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1321_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1609_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1624_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1610_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1611_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg988_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1534_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1584_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1626_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1598_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1612_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg969_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1536_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg990_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg998_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1650_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1484_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1539_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1002_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1592_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg401_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1589_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1488_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1649_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg405_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg375_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1491_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1545_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1602_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1637_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1493_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg166_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1495_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1548_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1549_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1614_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1629_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg409_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1577_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1505_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1010_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1529_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1579_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1642_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1329_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1433_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1558_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No126_out);

SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1321_out;
SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1322_out;
SharedReg1643_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1643_out;
SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg941_out;
SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg943_out;
SharedReg128_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg128_out;
SharedReg1644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1557_out;
SharedReg1328_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1328_out;
SharedReg1559_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1559_out;
SharedReg1435_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1435_out;
SharedReg1618_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1618_out;
SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg943_out;
SharedReg944_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg944_out;
SharedReg1324_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1324_out;
SharedReg1620_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1620_out;
SharedReg173_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg173_out;
SharedReg1019_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1019_out;
SharedReg947_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg947_out;
SharedReg1622_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1623_out;
SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1322_out;
SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1321_out;
SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1322_out;
SharedReg1326_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1326_out;
SharedReg1582_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1582_out;
SharedReg177_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg177_out;
SharedReg1341_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1341_out;
SharedReg968_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg968_out;
SharedReg969_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg969_out;
SharedReg1627_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1627_out;
SharedReg989_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg989_out;
SharedReg1587_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1537_out;
SharedReg998_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg998_out;
SharedReg1538_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1538_out;
SharedReg396_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg396_out;
SharedReg155_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg155_out;
SharedReg1651_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1540_out;
SharedReg972_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg972_out;
SharedReg1006_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1006_out;
SharedReg1001_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1001_out;
SharedReg1002_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1002_out;
SharedReg1543_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1544_out;
SharedReg980_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg980_out;
SharedReg164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg164_out;
SharedReg979_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg979_out;
SharedReg410_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg410_out;
SharedReg1546_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1546_out;
SharedReg166_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg166_out;
SharedReg411_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg411_out;
SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg167_out;
SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1011_out;
SharedReg1575_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1576_out;
SharedReg168_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg168_out;
SharedReg1578_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1578_out;
SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1011_out;
SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg167_out;
SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg940_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1559_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1435_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1618_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg944_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1324_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1620_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg173_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1019_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg947_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1643_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1622_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1623_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1321_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1322_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1326_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1582_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg177_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1341_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg968_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg969_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1627_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg989_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1587_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1537_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg998_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1538_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg396_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg155_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1651_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg941_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1540_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg972_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1006_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1001_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1002_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1543_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1544_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg980_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg979_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg943_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg410_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1546_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg166_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg411_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1575_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1576_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg168_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg128_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1578_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1011_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg167_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg940_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1557_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1328_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product32_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_5_impl_out,
                 X => Delay1No128_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg439_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg439_out;
SharedReg1387_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1387_out;
SharedReg1577_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1577_out;
SharedReg1038_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1038_out;
SharedReg1529_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1590_out;
SharedReg968_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg968_out;
SharedReg1598_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1505_out;
SharedReg1006_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1006_out;
SharedReg1326_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1326_out;
SharedReg1558_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1558_out;
SharedReg162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg162_out;
SharedReg1645_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1645_out;
SharedReg974_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg974_out;
SharedReg1619_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1607_out;
SharedReg1002_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1002_out;
SharedReg1530_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1608_out;
SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg998_out;
SharedReg1609_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1611_out;
SharedReg1020_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1020_out;
SharedReg1534_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1612_out;
SharedReg1028_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1028_out;
SharedReg1536_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1536_out;
SharedReg1022_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1022_out;
SharedReg1373_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1373_out;
SharedReg1650_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1650_out;
SharedReg183_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg183_out;
SharedReg1484_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1539_out;
SharedReg1377_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1377_out;
SharedReg431_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg431_out;
SharedReg1589_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1647_out;
SharedReg435_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg435_out;
SharedReg403_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg403_out;
SharedReg1491_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1493_out;
SharedReg194_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg194_out;
SharedReg1495_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1629_out;
   MUX_Product32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg439_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1387_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1598_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1592_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1637_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1505_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1006_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1326_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1558_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1645_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg974_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1577_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1619_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1606_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1607_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1002_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1530_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1580_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1608_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg998_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1609_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1038_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1624_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1610_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1611_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1020_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1534_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1584_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1626_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1612_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1028_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1536_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1529_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1022_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1373_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1650_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg183_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1484_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1539_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1377_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg431_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1589_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1488_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1579_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1649_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1647_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg435_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg403_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1491_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1545_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1602_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1493_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg194_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1495_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1642_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1548_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1549_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1614_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1629_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1596_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1590_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg968_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_5_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_0_out,
                 Y => Delay1No128_out);

SharedReg1575_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1576_out;
SharedReg197_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg197_out;
SharedReg1578_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1578_out;
SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1039_out;
SharedReg409_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg968_out;
SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg998_out;
SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg999_out;
SharedReg1643_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1643_out;
SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg968_out;
SharedReg969_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg969_out;
SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg971_out;
SharedReg158_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg158_out;
SharedReg1644_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1557_out;
SharedReg1005_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1005_out;
SharedReg1559_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1559_out;
SharedReg1328_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1328_out;
SharedReg1618_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1618_out;
SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg971_out;
SharedReg972_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg972_out;
SharedReg1001_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1001_out;
SharedReg1620_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1620_out;
SharedReg416_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg416_out;
SharedReg1047_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1047_out;
SharedReg975_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg975_out;
SharedReg1622_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1623_out;
SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg999_out;
SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg998_out;
SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg999_out;
SharedReg1003_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1003_out;
SharedReg1582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1582_out;
SharedReg420_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg420_out;
SharedReg989_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg989_out;
SharedReg1027_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1028_out;
SharedReg1627_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1627_out;
SharedReg1021_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1021_out;
SharedReg1587_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1537_out;
SharedReg1373_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1373_out;
SharedReg1538_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1538_out;
SharedReg426_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg426_out;
SharedReg184_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg184_out;
SharedReg1651_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1540_out;
SharedReg1031_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1031_out;
SharedReg1381_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1381_out;
SharedReg1376_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1376_out;
SharedReg1377_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1377_out;
SharedReg1543_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1544_out;
SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1039_out;
SharedReg192_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg192_out;
SharedReg1037_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1037_out;
SharedReg440_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg440_out;
SharedReg1546_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1546_out;
SharedReg194_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg194_out;
SharedReg441_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg441_out;
SharedReg195_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg195_out;
SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1386_out;
SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1386_out;
   MUX_Product32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1575_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1576_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg969_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg158_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1644_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1557_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1005_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1559_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1328_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1618_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg197_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg971_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg972_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1001_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1620_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg416_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1047_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg975_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1622_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1623_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1578_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1003_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg420_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg989_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1027_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1028_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1627_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1021_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1587_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1537_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1373_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1538_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg426_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg184_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1651_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1540_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1031_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1381_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg409_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1376_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1377_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1543_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1544_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1039_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg192_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1037_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg440_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1546_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg194_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg968_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg441_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg195_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1386_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg999_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1643_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_5_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product32_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_6_impl_out,
                 X => Delay1No130_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1493_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1493_out;
SharedReg221_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg1495_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1629_out;
SharedReg222_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg222_out;
SharedReg1070_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1070_out;
SharedReg1577_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1577_out;
SharedReg1385_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1385_out;
SharedReg1529_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1590_out;
SharedReg1027_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1027_out;
SharedReg1598_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1505_out;
SharedReg1381_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1381_out;
SharedReg1003_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1003_out;
SharedReg1558_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1558_out;
SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg191_out;
SharedReg1645_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1645_out;
SharedReg1032_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1032_out;
SharedReg1619_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1607_out;
SharedReg1377_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1377_out;
SharedReg1530_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1608_out;
SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1373_out;
SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1373_out;
SharedReg1609_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1611_out;
SharedReg1048_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1048_out;
SharedReg1534_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1612_out;
SharedReg1058_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1058_out;
SharedReg1536_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1536_out;
SharedReg1395_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1395_out;
SharedReg1295_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1295_out;
SharedReg1650_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1650_out;
SharedReg210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg210_out;
SharedReg1484_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1539_out;
SharedReg1299_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1299_out;
SharedReg240_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg240_out;
SharedReg1589_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1647_out;
SharedReg244_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg244_out;
SharedReg433_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg433_out;
SharedReg1491_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1602_out;
   MUX_Product32_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1493_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1385_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1529_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1579_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1642_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1596_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1590_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1027_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1598_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1592_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1637_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1495_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1505_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1381_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1003_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1558_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1645_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1032_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1619_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1606_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1607_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1548_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1377_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1530_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1580_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1608_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1373_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1609_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1624_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1610_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1611_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1549_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1048_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1534_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1584_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1626_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1612_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1058_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1536_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1395_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1295_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1650_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1614_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1484_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1539_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1299_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg240_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1589_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1488_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1649_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1647_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg244_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1629_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg433_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1491_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1545_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1602_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg222_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1070_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1577_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_6_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_0_out,
                 Y => Delay1No130_out);

SharedReg249_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg1546_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1546_out;
SharedReg438_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg438_out;
SharedReg250_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg250_out;
SharedReg439_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg439_out;
SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1069_out;
SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1069_out;
SharedReg1575_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1576_out;
SharedReg441_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg441_out;
SharedReg1578_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1578_out;
SharedReg1386_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1386_out;
SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg195_out;
SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1027_out;
SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1373_out;
SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1374_out;
SharedReg1643_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1643_out;
SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1028_out;
SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1030_out;
SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg187_out;
SharedReg1644_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1557_out;
SharedReg1380_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1380_out;
SharedReg1559_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1559_out;
SharedReg1005_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1005_out;
SharedReg1618_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1618_out;
SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1031_out;
SharedReg1376_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1376_out;
SharedReg1620_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1620_out;
SharedReg202_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg202_out;
SharedReg1393_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1393_out;
SharedReg1033_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1033_out;
SharedReg1622_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1623_out;
SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1374_out;
SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1373_out;
SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1374_out;
SharedReg1378_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1378_out;
SharedReg1582_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1582_out;
SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg204_out;
SharedReg1021_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1021_out;
SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1057_out;
SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1058_out;
SharedReg1627_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1627_out;
SharedReg1394_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1394_out;
SharedReg1587_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1537_out;
SharedReg1295_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1295_out;
SharedReg1538_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1538_out;
SharedReg235_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg235_out;
SharedReg211_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg211_out;
SharedReg1651_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1540_out;
SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1061_out;
SharedReg1303_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1303_out;
SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1060_out;
SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1061_out;
SharedReg1543_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1544_out;
SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1069_out;
SharedReg219_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg219_out;
SharedReg1067_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1067_out;
   MUX_Product32_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1546_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1578_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1386_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1643_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1027_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1028_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg438_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1644_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1557_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1380_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1559_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1005_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1618_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1030_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1031_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1376_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg250_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1620_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg202_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1393_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1033_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1622_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1623_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1373_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1378_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg439_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1582_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1021_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1627_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1394_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1587_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1537_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1295_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1538_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg235_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg211_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1651_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1540_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1303_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1061_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1543_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1544_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1069_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg219_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1067_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1575_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1576_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg441_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_6_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product32_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_7_impl_out,
                 X => Delay1No132_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1649_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1647_out;
SharedReg270_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg270_out;
SharedReg217_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg217_out;
SharedReg1491_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1493_out;
SharedReg247_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg247_out;
SharedReg1495_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1629_out;
SharedReg248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg248_out;
SharedReg1309_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1309_out;
SharedReg1577_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1577_out;
SharedReg1307_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1307_out;
SharedReg1529_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1590_out;
SharedReg1057_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1057_out;
SharedReg1598_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1505_out;
SharedReg1303_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1303_out;
SharedReg1378_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1378_out;
SharedReg1558_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1558_out;
SharedReg218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg218_out;
SharedReg1645_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1645_out;
SharedReg1062_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1062_out;
SharedReg1619_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1607_out;
SharedReg1299_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1299_out;
SharedReg1530_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1608_out;
SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1295_out;
SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1295_out;
SharedReg1609_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1611_out;
SharedReg1077_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1077_out;
SharedReg1534_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1612_out;
SharedReg1087_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1087_out;
SharedReg1536_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1536_out;
SharedReg1315_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1315_out;
SharedReg1086_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1086_out;
SharedReg1650_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1650_out;
SharedReg235_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg235_out;
SharedReg1484_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1539_out;
SharedReg1090_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1090_out;
SharedReg266_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg266_out;
SharedReg1589_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1488_out;
   MUX_Product32_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1649_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1647_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1548_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1549_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1614_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1629_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1309_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1577_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1307_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1529_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1579_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg270_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1642_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1596_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1590_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1057_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1598_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1592_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1637_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1505_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1303_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1378_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg217_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1558_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1645_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1062_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1619_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1606_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1607_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1299_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1530_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1580_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1491_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1608_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1295_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1609_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1624_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1610_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1611_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1077_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1534_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1584_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1545_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1626_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1612_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1087_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1536_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1315_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1086_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1650_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg235_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1484_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1539_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1602_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1090_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg266_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1589_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1488_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1493_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg247_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1495_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_7_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_7_impl_0_out,
                 Y => Delay1No132_out);

SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1298_out;
SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1299_out;
SharedReg1543_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1544_out;
SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1308_out;
SharedReg245_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg245_out;
SharedReg1306_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg275_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg275_out;
SharedReg1546_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1546_out;
SharedReg221_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg221_out;
SharedReg276_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg276_out;
SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg222_out;
SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1308_out;
SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1308_out;
SharedReg1575_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1576_out;
SharedReg223_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg223_out;
SharedReg1578_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1578_out;
SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1308_out;
SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg222_out;
SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1057_out;
SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1295_out;
SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1296_out;
SharedReg1643_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1643_out;
SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1057_out;
SharedReg1058_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1058_out;
SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1060_out;
SharedReg214_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg214_out;
SharedReg1644_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1557_out;
SharedReg1302_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1302_out;
SharedReg1559_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1559_out;
SharedReg1380_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1380_out;
SharedReg1618_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1618_out;
SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1060_out;
SharedReg1061_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1061_out;
SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1298_out;
SharedReg1620_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1620_out;
SharedReg227_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg227_out;
SharedReg1313_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1313_out;
SharedReg1063_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1063_out;
SharedReg1622_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1623_out;
SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1296_out;
SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1295_out;
SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1296_out;
SharedReg1300_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1300_out;
SharedReg1582_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1582_out;
SharedReg229_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg229_out;
SharedReg1394_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1394_out;
SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1086_out;
SharedReg1087_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1087_out;
SharedReg1627_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1627_out;
SharedReg1314_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1314_out;
SharedReg1587_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1537_out;
SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1086_out;
SharedReg1538_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1538_out;
SharedReg261_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg261_out;
SharedReg236_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_60_cast <= SharedReg236_out;
SharedReg1651_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1540_out;
SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1299_out;
SharedReg1094_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1094_out;
   MUX_Product32_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1575_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1576_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg223_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1578_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg222_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1543_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1643_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1057_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1058_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg214_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1644_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1557_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1544_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1302_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1559_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1380_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1618_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1060_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1061_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1298_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1620_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg227_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1313_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1308_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1063_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1622_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1623_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1295_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1296_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1300_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1582_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg229_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1394_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg245_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1087_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1627_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1314_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1587_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1537_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1086_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1538_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg261_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg236_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1651_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1540_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1299_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1094_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg275_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1546_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg221_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_7_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_7_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product32_8_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product32_8_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product32_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_8_impl_out,
                 X => Delay1No134_out_to_Product32_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product32_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1650_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1650_out;
SharedReg261_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg261_out;
SharedReg1484_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1484_out;
SharedReg1539_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1539_out;
SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1461_out;
SharedReg461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg461_out;
SharedReg1589_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1589_out;
SharedReg1488_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1488_out;
SharedReg1649_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1649_out;
SharedReg1647_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1647_out;
SharedReg465_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg465_out;
SharedReg242_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg242_out;
SharedReg1491_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1491_out;
SharedReg1545_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1545_out;
SharedReg1602_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1602_out;
SharedReg1493_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1493_out;
SharedReg273_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg273_out;
SharedReg1495_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1495_out;
SharedReg1548_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1548_out;
SharedReg1549_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1549_out;
SharedReg1614_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1614_out;
SharedReg1629_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1629_out;
SharedReg469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg469_out;
SharedReg1469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1469_out;
SharedReg1577_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1577_out;
SharedReg1467_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1467_out;
SharedReg1529_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1529_out;
SharedReg1579_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1579_out;
SharedReg1642_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1642_out;
SharedReg1596_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1596_out;
SharedReg1590_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1590_out;
SharedReg1295_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1295_out;
SharedReg1598_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1598_out;
SharedReg1592_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1592_out;
SharedReg1637_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1637_out;
SharedReg1505_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1505_out;
SharedReg1463_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1463_out;
SharedReg1300_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1300_out;
SharedReg1558_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1558_out;
SharedReg269_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg269_out;
SharedReg1645_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1645_out;
SharedReg1092_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1092_out;
SharedReg1619_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1619_out;
SharedReg1606_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1606_out;
SharedReg1607_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1607_out;
SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1461_out;
SharedReg1530_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1530_out;
SharedReg1580_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1580_out;
SharedReg1608_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1608_out;
SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1457_out;
SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1457_out;
SharedReg1609_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1609_out;
SharedReg1624_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1624_out;
SharedReg1610_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1610_out;
SharedReg1611_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1611_out;
SharedReg1106_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1106_out;
SharedReg1534_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1534_out;
SharedReg1584_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1584_out;
SharedReg1626_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1626_out;
SharedReg1612_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1612_out;
SharedReg1458_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1458_out;
SharedReg1536_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1536_out;
SharedReg1477_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1477_out;
SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1457_out;
   MUX_Product32_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1650_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg261_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg465_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg242_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1491_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1545_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1602_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1493_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg273_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1495_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1548_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1549_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1484_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1614_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1629_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1469_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1577_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1467_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1529_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1579_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1642_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1596_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1539_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1590_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1295_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1598_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1592_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1637_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1505_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1463_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1300_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1558_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg269_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1645_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1092_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1619_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1606_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1607_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1530_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1580_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1608_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg461_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1609_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1624_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1610_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1611_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1106_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1534_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1584_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1626_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1612_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1589_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1458_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1536_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1477_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1457_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1488_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1649_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1647_out_to_MUX_Product32_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_8_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_8_impl_0_out,
                 Y => Delay1No134_out);

SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1457_out;
SharedReg1538_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1538_out;
SharedReg457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg457_out;
SharedReg262_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg1651_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1651_out;
SharedReg1540_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1540_out;
SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1090_out;
SharedReg1463_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1463_out;
SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1460_out;
SharedReg1461_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1461_out;
SharedReg1543_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1543_out;
SharedReg1544_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1544_out;
SharedReg1099_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1099_out;
SharedReg245_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg245_out;
SharedReg1306_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1306_out;
SharedReg470_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg470_out;
SharedReg1546_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1546_out;
SharedReg273_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg273_out;
SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg276_out;
SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg274_out;
SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1468_out;
SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1468_out;
SharedReg1575_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1575_out;
SharedReg1576_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1576_out;
SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg276_out;
SharedReg1578_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1578_out;
SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1468_out;
SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg274_out;
SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1086_out;
SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1457_out;
SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1458_out;
SharedReg1643_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1643_out;
SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1086_out;
SharedReg1087_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1087_out;
SharedReg1298_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1298_out;
SharedReg265_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg265_out;
SharedReg1644_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1644_out;
SharedReg1557_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1557_out;
SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1093_out;
SharedReg1559_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1559_out;
SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1093_out;
SharedReg1618_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1618_out;
SharedReg1089_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1090_out;
SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1460_out;
SharedReg1620_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1620_out;
SharedReg280_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg280_out;
SharedReg1475_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1475_out;
SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1093_out;
SharedReg1622_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1622_out;
SharedReg1623_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1623_out;
SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1458_out;
SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1457_out;
SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1458_out;
SharedReg1462_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1462_out;
SharedReg1582_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1582_out;
SharedReg479_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg479_out;
SharedReg1107_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1107_out;
SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1457_out;
SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1458_out;
SharedReg1627_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1627_out;
SharedReg1476_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1476_out;
SharedReg1587_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1587_out;
SharedReg1537_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1537_out;
   MUX_Product32_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1538_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1543_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1544_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1099_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg245_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1306_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg470_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1546_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg273_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1575_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1576_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg276_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1578_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1468_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg274_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg262_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1643_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1086_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1087_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1298_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg265_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1644_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1557_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1559_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1651_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1618_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1089_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1620_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg280_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1475_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1093_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1622_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1540_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1623_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1462_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1582_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg479_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1107_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1457_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1458_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1090_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1627_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1476_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1587_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1537_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1463_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1460_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1461_out_to_MUX_Product32_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_8_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_8_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Subtract3_8_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Subtract3_8_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Subtract3_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_8_impl_out,
                 X => Delay1No136_out_to_Subtract3_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Subtract3_8_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1058_out;
SharedReg1057_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1057_out;
SharedReg1296_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1296_out;
SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg1289_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1289_out;
SharedReg848_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg848_out;
SharedReg214_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg214_out;
SharedReg1255_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1255_out;
SharedReg1060_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1060_out;
SharedReg447_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg447_out;
SharedReg813_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg813_out;
SharedReg652_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg652_out;
SharedReg1275_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1275_out;
SharedReg241_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg241_out;
SharedReg210_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg210_out;
SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1067_out;
SharedReg247_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg247_out;
SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1067_out;
SharedReg658_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg658_out;
SharedReg1290_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1290_out;
SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg817_out;
SharedReg1304_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1304_out;
SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg821_out;
SharedReg244_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg244_out;
SharedReg1064_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1064_out;
SharedReg457_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg457_out;
SharedReg468_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg468_out;
SharedReg226_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg226_out;
SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1058_out;
SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg237_out;
SharedReg212_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg212_out;
SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg821_out;
SharedReg1303_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1303_out;
SharedReg653_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg653_out;
SharedReg633_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg633_out;
SharedReg240_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg240_out;
SharedReg431_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg431_out;
SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1380_out;
SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1380_out;
SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg817_out;
SharedReg636_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg636_out;
SharedReg1235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1235_out;
SharedReg1_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg11_out;
SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_49_cast <= SharedReg631_out;
SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_50_cast <= SharedReg631_out;
SharedReg_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_51_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_52_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_53_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_54_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_55_cast <= SharedReg7_out;
SharedReg12_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_56_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_57_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_58_cast <= SharedReg13_out;
SharedReg252_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_59_cast <= SharedReg252_out;
SharedReg1075_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1075_out;
SharedReg272_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_61_cast <= SharedReg272_out;
SharedReg826_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_62_cast <= SharedReg826_out;
SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_63_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_64_cast <= SharedReg10_out;
   MUX_Subtract3_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg447_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg813_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg652_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1275_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg241_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg210_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg247_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1067_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg658_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1057_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1290_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1304_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg244_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1064_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg457_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg468_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg226_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1058_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1296_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg212_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg821_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1303_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg653_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg633_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg240_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg431_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1380_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg237_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg817_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg636_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1235_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg3_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg17_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg6_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg11_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg631_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1289_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg2_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg14_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg4_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg12_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg16_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg13_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg252_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1075_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg848_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg272_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg826_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg7_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg10_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg214_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1255_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1060_out_to_MUX_Subtract3_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract3_8_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_8_impl_0_out,
                 Y => Delay1No136_out);

SharedReg277_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg1101_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1101_out;
SharedReg1320_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1320_out;
SharedReg1113_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg287_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg287_out;
Delay43No17_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_6_cast <= Delay43No17_out;
SharedReg664_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg664_out;
SharedReg233_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg233_out;
SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1266_out;
SharedReg1319_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1319_out;
SharedReg218_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg218_out;
SharedReg1260_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1260_out;
SharedReg1278_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1278_out;
SharedReg660_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg660_out;
SharedReg236_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg236_out;
SharedReg241_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg241_out;
SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1057_out;
SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg210_out;
SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1057_out;
SharedReg652_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg652_out;
SharedReg847_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg847_out;
SharedReg1273_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1273_out;
SharedReg1065_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1065_out;
SharedReg828_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg828_out;
SharedReg234_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg234_out;
SharedReg1082_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1082_out;
SharedReg459_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg459_out;
SharedReg261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg261_out;
SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg210_out;
SharedReg1109_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1109_out;
SharedReg284_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg284_out;
SharedReg254_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg254_out;
SharedReg1255_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1255_out;
SharedReg1114_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1114_out;
SharedReg833_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg833_out;
SharedReg813_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg813_out;
SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg235_out;
SharedReg1058_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1058_out;
SharedReg1297_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1297_out;
SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1266_out;
SharedReg1261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1261_out;
SharedReg1238_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1238_out;
SharedReg19_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg29_out;
SharedReg815_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_49_cast <= SharedReg815_out;
SharedReg1259_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1259_out;
SharedReg18_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_51_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_52_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_53_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_54_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_55_cast <= SharedReg25_out;
SharedReg30_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_56_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_57_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_58_cast <= SharedReg31_out;
SharedReg221_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_59_cast <= SharedReg221_out;
SharedReg1308_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1308_out;
SharedReg274_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_61_cast <= SharedReg274_out;
Delay41No25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_62_cast <= Delay41No25_out;
SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_63_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_64_cast <= SharedReg28_out;
   MUX_Subtract3_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1101_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg218_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1260_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1278_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg660_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg236_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg241_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1057_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg652_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1320_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg847_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1273_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1065_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg828_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg234_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1082_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg459_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg210_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1109_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg284_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg254_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1255_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1114_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg833_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg813_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg235_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1058_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1297_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg287_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1261_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1238_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg19_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg21_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg35_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg24_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg29_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg815_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1259_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => Delay43No17_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg18_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg20_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg32_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg22_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg30_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg34_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg31_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg221_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1308_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg664_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg274_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => Delay41No25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg25_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg28_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg233_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1266_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1319_out_to_MUX_Subtract3_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract3_8_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_8_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Subtract5_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_4_impl_out,
                 X => Delay1No138_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg757_out;
SharedReg977_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg977_out;
SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg761_out;
SharedReg163_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg163_out;
SharedReg1329_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1329_out;
SharedReg194_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg194_out;
SharedReg1323_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1323_out;
SharedReg172_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg172_out;
SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg941_out;
SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg370_out;
SharedReg126_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg126_out;
SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg761_out;
SharedReg590_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg590_out;
SharedReg1216_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1216_out;
SharedReg570_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg570_out;
SharedReg373_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg373_out;
SharedReg129_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg129_out;
SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1435_out;
SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1435_out;
SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg757_out;
SharedReg573_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg573_out;
SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1175_out;
SharedReg1_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg13_out;
SharedReg359_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg359_out;
SharedReg927_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg927_out;
SharedReg134_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg134_out;
SharedReg746_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg746_out;
SharedReg1188_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1188_out;
SharedReg556_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg556_out;
SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg368_out;
SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg941_out;
SharedReg940_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg940_out;
SharedReg1322_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1322_out;
SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg370_out;
SharedReg360_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg360_out;
SharedReg929_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg929_out;
SharedReg128_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg128_out;
SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1175_out;
SharedReg943_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg943_out;
SharedReg115_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg115_out;
SharedReg733_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg733_out;
SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1195_out;
SharedReg1338_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1338_out;
SharedReg1001_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1001_out;
SharedReg569_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg569_out;
SharedReg401_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg401_out;
SharedReg568_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg568_out;
SharedReg574_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg574_out;
SharedReg585_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg585_out;
SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1195_out;
SharedReg402_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg402_out;
SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg368_out;
SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg979_out;
SharedReg408_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg408_out;
SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg979_out;
SharedReg1230_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1230_out;
SharedReg777_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg777_out;
   MUX_Subtract5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg977_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg126_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg590_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1216_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg570_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg373_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg129_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1435_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg757_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg761_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg573_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg3_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg17_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg6_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg11_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg12_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg16_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg13_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg163_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg359_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg927_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg134_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg746_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1188_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg556_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg940_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1322_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1329_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg360_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg929_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg128_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1175_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg943_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg115_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg733_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1338_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg194_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1001_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg569_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg401_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg568_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg574_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg585_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1195_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg402_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg368_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1323_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg408_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg979_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1230_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg777_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg172_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg941_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg370_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract5_4_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_0_out,
                 Y => Delay1No138_out);

SharedReg1213_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1213_out;
SharedReg1330_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1330_out;
SharedReg768_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg768_out;
SharedReg182_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg964_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg964_out;
SharedReg154_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg1002_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1002_out;
SharedReg124_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg124_out;
SharedReg992_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg992_out;
SharedReg180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg180_out;
SharedReg416_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg416_out;
SharedReg1195_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1195_out;
SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg773_out;
SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg773_out;
SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg753_out;
SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg368_out;
SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg368_out;
SharedReg941_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg941_out;
SharedReg1323_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1323_out;
SharedReg1206_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1206_out;
SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1201_out;
SharedReg1178_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1178_out;
SharedReg19_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg31_out;
SharedReg355_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg355_out;
SharedReg1441_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1441_out;
SharedReg136_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg136_out;
Delay41No21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_34_cast <= Delay41No21_out;
SharedReg1191_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1191_out;
SharedReg745_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg745_out;
SharedReg138_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg138_out;
SharedReg954_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg954_out;
SharedReg966_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg966_out;
SharedReg1346_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1346_out;
SharedReg395_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg395_out;
SharedReg345_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg345_out;
SharedReg1324_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1324_out;
SharedReg121_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg121_out;
SharedReg1186_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1186_out;
SharedReg1452_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1452_out;
SharedReg132_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg132_out;
SharedReg1180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1180_out;
SharedReg576_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg576_out;
SharedReg971_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg971_out;
SharedReg963_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg963_out;
SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg753_out;
SharedReg392_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg392_out;
SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg569_out;
SharedReg568_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg568_out;
SharedReg1208_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1208_out;
SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1201_out;
SharedReg155_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg155_out;
SharedReg402_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg402_out;
SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1321_out;
SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg368_out;
SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1321_out;
SharedReg787_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg787_out;
SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg773_out;
   MUX_Subtract5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1213_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1330_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg416_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1195_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg941_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1323_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1206_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg768_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1178_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg19_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg35_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg24_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg29_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg30_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg34_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg182_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg355_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1441_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg136_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay41No21_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1191_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg745_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg138_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg954_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg966_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1346_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg964_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg395_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg345_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1324_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg121_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1186_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1452_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg132_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg576_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg971_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg154_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg963_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg753_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg392_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg568_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1208_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1201_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg155_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg402_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1002_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg368_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1321_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg787_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg773_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg124_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg992_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg180_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract5_4_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Subtract8_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_2_impl_out,
                 X => Delay1No140_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast);

SharedReg528_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg528_out;
SharedReg100_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg322_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg322_out;
SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg889_out;
SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg889_out;
SharedReg717_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg717_out;
SharedReg531_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg531_out;
SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1135_out;
SharedReg1_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg13_out;
SharedReg84_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg84_out;
SharedReg1417_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1417_out;
SharedReg76_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg76_out;
SharedReg706_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg706_out;
SharedReg1148_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1148_out;
SharedReg514_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg514_out;
SharedReg317_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg317_out;
SharedReg883_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg883_out;
SharedReg882_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg882_out;
SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1348_out;
SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg319_out;
SharedReg307_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg307_out;
SharedReg1419_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1419_out;
SharedReg321_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg321_out;
SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1135_out;
SharedReg885_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg885_out;
SharedReg310_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg310_out;
SharedReg693_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg693_out;
SharedReg522_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg522_out;
SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1135_out;
SharedReg323_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg323_out;
SharedReg66_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg66_out;
SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg893_out;
SharedReg329_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg329_out;
SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg893_out;
SharedReg892_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg892_out;
SharedReg331_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg331_out;
SharedReg697_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg697_out;
SharedReg1356_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1356_out;
SharedReg701_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg701_out;
SharedReg326_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg326_out;
SharedReg1355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1355_out;
SharedReg355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg355_out;
SharedReg912_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg912_out;
SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg529_out;
SharedReg111_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg111_out;
SharedReg716_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg716_out;
SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg529_out;
SharedReg918_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg918_out;
SharedReg925_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg925_out;
SharedReg105_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg105_out;
SharedReg112_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg112_out;
SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1348_out;
SharedReg97_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg97_out;
SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg319_out;
SharedReg721_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg721_out;
SharedReg548_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg548_out;
SharedReg1176_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1176_out;
   MUX_Subtract8_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg528_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg6_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg16_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg84_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1417_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg76_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg706_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg322_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1148_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg514_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg317_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg883_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg882_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg307_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1419_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg321_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg885_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg310_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg693_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg522_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg323_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg66_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg329_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg889_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg893_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg892_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg331_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg697_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1356_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg701_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg326_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg355_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg912_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg717_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg111_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg716_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg529_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg918_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg925_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg105_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg112_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1348_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg97_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg531_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg319_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg721_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg548_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1176_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1135_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg3_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract8_2_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_2_impl_0_out,
                 Y => Delay1No140_out);

SharedReg713_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg713_out;
SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg883_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg1349_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1349_out;
SharedReg1166_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1166_out;
SharedReg1161_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1161_out;
SharedReg1138_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1138_out;
SharedReg19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg31_out;
SharedReg302_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg302_out;
SharedReg1413_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1413_out;
SharedReg78_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg78_out;
Delay41No19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_20_cast <= Delay41No19_out;
SharedReg1151_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1151_out;
SharedReg705_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg705_out;
SharedReg80_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg80_out;
SharedReg896_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg896_out;
SharedReg908_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg908_out;
SharedReg1372_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1372_out;
SharedReg342_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg342_out;
SharedReg68_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg68_out;
SharedReg1350_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1350_out;
SharedReg93_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg93_out;
SharedReg1146_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1146_out;
SharedReg1371_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1371_out;
SharedReg74_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg74_out;
SharedReg1140_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1140_out;
SharedReg1148_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1148_out;
SharedReg1141_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1141_out;
SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg318_out;
SharedReg323_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg323_out;
SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg882_out;
SharedReg66_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg66_out;
SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1347_out;
SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg882_out;
SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg318_out;
SharedReg1153_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1153_out;
SharedReg891_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg891_out;
SharedReg708_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg708_out;
SharedReg94_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg94_out;
SharedReg906_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg906_out;
SharedReg95_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg95_out;
SharedReg1432_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1432_out;
SharedReg541_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg541_out;
SharedReg343_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg343_out;
SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1160_out;
SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1160_out;
SharedReg939_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg939_out;
SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1347_out;
SharedReg365_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg365_out;
SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg317_out;
SharedReg932_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg932_out;
SharedReg119_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg119_out;
SharedReg361_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg361_out;
SharedReg1155_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1155_out;
SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg733_out;
SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg733_out;
   MUX_Subtract8_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg713_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg35_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg34_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg31_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg302_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1413_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg78_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay41No19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1151_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg705_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg80_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg896_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg908_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1372_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg342_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg68_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1350_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg93_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg883_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1146_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1371_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg74_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1140_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1148_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1141_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg323_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg66_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1349_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg882_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg318_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1153_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg891_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg708_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg94_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg906_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg95_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1432_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1166_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg541_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg343_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1160_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg939_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1347_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg365_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg317_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg932_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg119_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1161_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg361_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1155_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg733_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1138_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg19_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg21_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract8_2_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_2_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract9_7_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract9_7_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract9_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_7_impl_out,
                 X => Delay1No142_out_to_Subtract9_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract9_7_impl_parent_implementedSystem_port_1_cast);

SharedReg430_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg430_out;
SharedReg1235_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1235_out;
SharedReg1030_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1030_out;
SharedReg418_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg418_out;
SharedReg793_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg793_out;
SharedReg1255_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1255_out;
SharedReg1312_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1312_out;
SharedReg432_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg432_out;
SharedReg183_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg183_out;
SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1037_out;
SharedReg438_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg438_out;
SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1037_out;
SharedReg1270_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1270_out;
SharedReg817_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg817_out;
SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg797_out;
SharedReg1382_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1382_out;
SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg801_out;
SharedReg435_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg435_out;
SharedReg1034_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1034_out;
SharedReg247_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg247_out;
SharedReg1375_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1375_out;
SharedReg201_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg201_out;
SharedReg1028_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1028_out;
SharedReg428_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg428_out;
SharedReg185_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg185_out;
SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg801_out;
SharedReg632_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg632_out;
SharedReg1256_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1256_out;
SharedReg612_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_29_cast <= SharedReg612_out;
SharedReg431_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_30_cast <= SharedReg431_out;
SharedReg188_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_31_cast <= SharedReg188_out;
SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1005_out;
SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1005_out;
SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_34_cast <= SharedReg797_out;
SharedReg615_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_35_cast <= SharedReg615_out;
SharedReg1215_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1215_out;
SharedReg1_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_38_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_39_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_40_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_41_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_42_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_43_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_44_cast <= SharedReg13_out;
SharedReg414_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_45_cast <= SharedReg414_out;
SharedReg985_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_46_cast <= SharedReg985_out;
SharedReg193_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_47_cast <= SharedReg193_out;
SharedReg786_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_48_cast <= SharedReg786_out;
SharedReg10_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_49_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_50_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_51_cast <= SharedReg8_out;
SharedReg614_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_52_cast <= SharedReg614_out;
SharedReg622_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_53_cast <= SharedReg622_out;
SharedReg1067_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1067_out;
SharedReg1249_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1249_out;
SharedReg1248_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1248_out;
SharedReg619_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_57_cast <= SharedReg619_out;
SharedReg210_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_58_cast <= SharedReg210_out;
SharedReg1374_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1374_out;
SharedReg1373_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1373_out;
SharedReg1058_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1058_out;
SharedReg212_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_62_cast <= SharedReg212_out;
SharedReg828_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_63_cast <= SharedReg828_out;
SharedReg813_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_64_cast <= SharedReg813_out;
   MUX_Subtract9_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg430_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1235_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg438_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1270_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg817_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1382_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg435_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1034_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg247_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1030_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1375_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg201_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1028_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg428_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg185_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg801_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg632_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1256_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg612_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg431_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg418_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg188_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1005_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg797_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg615_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1215_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg3_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg17_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg6_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg793_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg11_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg12_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg16_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg13_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg414_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg985_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg193_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg786_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg10_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg9_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1255_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg8_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg614_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg622_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1067_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1249_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1248_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg619_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg210_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1374_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1373_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1312_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1058_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg212_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg828_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg813_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg432_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg183_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1037_out_to_MUX_Subtract9_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract9_7_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_7_impl_0_out,
                 Y => Delay1No142_out);

SharedReg208_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1246_out;
SharedReg1397_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1397_out;
SharedReg434_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg434_out;
SharedReg1240_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1240_out;
SharedReg639_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg639_out;
SharedReg1376_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1376_out;
SharedReg427_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg427_out;
SharedReg432_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg432_out;
SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1027_out;
SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg183_out;
SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1027_out;
SharedReg827_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg827_out;
SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg813_out;
SharedReg1253_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1253_out;
SharedReg1035_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1035_out;
SharedReg808_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg808_out;
SharedReg456_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg456_out;
SharedReg1053_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1053_out;
SharedReg210_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg210_out;
SharedReg1299_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1299_out;
SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg183_out;
SharedReg1080_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1080_out;
SharedReg232_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg232_out;
SharedReg227_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg227_out;
SharedReg1235_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1235_out;
SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg813_out;
SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg813_out;
SharedReg793_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_29_cast <= SharedReg793_out;
SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_30_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_31_cast <= SharedReg426_out;
SharedReg1028_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1028_out;
SharedReg1375_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1375_out;
SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1246_out;
SharedReg1241_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1241_out;
SharedReg1218_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1218_out;
SharedReg19_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_37_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_38_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_39_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_40_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_41_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_42_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_43_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_44_cast <= SharedReg31_out;
SharedReg166_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_45_cast <= SharedReg166_out;
SharedReg1011_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1011_out;
SharedReg195_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_47_cast <= SharedReg195_out;
Delay41No23_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_48_cast <= Delay41No23_out;
SharedReg28_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_49_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_50_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_51_cast <= SharedReg26_out;
SharedReg796_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_52_cast <= SharedReg796_out;
Delay37No42_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_53_cast <= Delay37No42_out;
SharedReg1069_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1069_out;
Delay43No15_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_55_cast <= Delay43No15_out;
SharedReg1251_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1251_out;
SharedReg805_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_57_cast <= SharedReg805_out;
SharedReg224_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_58_cast <= SharedReg224_out;
SharedReg1073_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1073_out;
SharedReg1084_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1084_out;
SharedReg1320_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1320_out;
SharedReg260_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_62_cast <= SharedReg260_out;
SharedReg643_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_63_cast <= SharedReg643_out;
SharedReg1257_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1257_out;
   MUX_Subtract9_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg827_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1253_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1035_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg808_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg456_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1053_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg210_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1397_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1299_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg183_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1080_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg232_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg227_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1235_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg813_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg793_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg434_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg426_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1028_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1375_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1246_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1241_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1218_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg19_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg21_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg35_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg24_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1240_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg29_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg30_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg34_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg31_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg166_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1011_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg195_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => Delay41No23_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg28_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg27_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg639_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg26_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg796_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => Delay37No42_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1069_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay43No15_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1251_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg805_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg224_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1073_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1084_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1376_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1320_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg260_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg643_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1257_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg427_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg432_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1027_out_to_MUX_Subtract9_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract9_7_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_7_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Subtract10_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_1_impl_out,
                 X => Delay1No144_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1115_out;
SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg306_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg306_out;
SharedReg870_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg870_out;
SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg686_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg686_out;
SharedReg1128_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1128_out;
SharedReg493_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg493_out;
SharedReg290_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg290_out;
SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg854_out;
SharedReg853_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg853_out;
SharedReg1401_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1401_out;
SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg292_out;
SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg54_out;
SharedReg873_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg873_out;
SharedReg294_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg294_out;
SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1115_out;
SharedReg856_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg856_out;
SharedReg57_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg57_out;
SharedReg673_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg673_out;
SharedReg501_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg501_out;
SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1115_out;
SharedReg296_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg296_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg36_out;
SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg864_out;
SharedReg302_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg302_out;
SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg864_out;
SharedReg863_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg863_out;
SharedReg304_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg304_out;
SharedReg677_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg677_out;
SharedReg1409_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1409_out;
SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg681_out;
SharedReg299_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg299_out;
SharedReg1408_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1408_out;
SharedReg868_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg868_out;
SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg53_out;
SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg854_out;
SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg292_out;
SharedReg38_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg38_out;
SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg681_out;
SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg506_out;
SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1136_out;
SharedReg898_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg898_out;
SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg506_out;
SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1136_out;
SharedReg884_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg884_out;
SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg505_out;
SharedReg321_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg321_out;
SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg505_out;
SharedReg507_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg507_out;
SharedReg322_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg322_out;
SharedReg71_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg71_out;
SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1407_out;
SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1407_out;
SharedReg697_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg697_out;
SharedReg510_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg510_out;
   MUX_Subtract10_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg870_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg686_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1128_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg493_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg290_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg853_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1401_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg873_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg294_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg856_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg57_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg673_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg501_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1115_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg296_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg36_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg302_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg864_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg863_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg304_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg677_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1409_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg299_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1408_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg868_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg46_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg53_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg854_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg292_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg38_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg681_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg898_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg506_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1136_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg884_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg321_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg505_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg507_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg322_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg71_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1407_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg697_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg510_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg306_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_1_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_1_impl_0_out,
                 Y => Delay1No144_out);

SharedReg1118_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1118_out;
SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg47_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg47_out;
SharedReg865_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg865_out;
SharedReg48_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg48_out;
Delay41No18_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast <= Delay41No18_out;
SharedReg1131_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1131_out;
SharedReg685_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg685_out;
SharedReg50_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg50_out;
SharedReg867_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg867_out;
SharedReg880_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg880_out;
SharedReg1427_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1427_out;
SharedReg316_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg316_out;
SharedReg38_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg38_out;
SharedReg1403_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1403_out;
SharedReg64_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg64_out;
SharedReg1126_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1126_out;
SharedReg1426_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1426_out;
SharedReg44_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg44_out;
SharedReg1120_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1120_out;
SharedReg1128_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1128_out;
SharedReg1121_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1121_out;
SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg291_out;
SharedReg296_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg296_out;
SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg853_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg1400_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1400_out;
SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg853_out;
SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg291_out;
SharedReg1133_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1133_out;
SharedReg862_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg862_out;
SharedReg688_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg688_out;
SharedReg65_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg65_out;
SharedReg878_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg878_out;
SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg853_out;
SharedReg314_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg314_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg36_out;
SharedReg876_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg876_out;
SharedReg62_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg62_out;
SharedReg308_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg308_out;
SharedReg1115_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1115_out;
SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg693_out;
SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg693_out;
SharedReg1347_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1347_out;
SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg693_out;
SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg693_out;
SharedReg904_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg904_out;
SharedReg694_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg694_out;
SharedReg92_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg92_out;
SharedReg1136_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1136_out;
SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg693_out;
SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg66_out;
SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg66_out;
SharedReg1401_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1401_out;
SharedReg884_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg884_out;
SharedReg1146_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1146_out;
SharedReg1141_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1141_out;
   MUX_Subtract10_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1118_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg865_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay41No18_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1131_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg685_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg50_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg867_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg880_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1427_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg316_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg38_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1403_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg64_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1126_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1426_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg44_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1120_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1128_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1121_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg296_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1400_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg291_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1133_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg862_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg688_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg65_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg878_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg853_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg314_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg876_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg62_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg308_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1115_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1347_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg904_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg694_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg92_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1136_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg693_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg66_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1401_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg884_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1146_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1141_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg47_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_1_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_1_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Subtract10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_3_impl_out,
                 X => Delay1No146_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg141_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg911_out;
SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg97_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg97_out;
SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg741_out;
SharedReg569_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg569_out;
SharedReg1196_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1196_out;
SharedReg549_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg549_out;
SharedReg348_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg348_out;
SharedReg100_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg100_out;
SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1354_out;
SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1354_out;
SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg737_out;
SharedReg552_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg552_out;
SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1155_out;
SharedReg1_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg13_out;
SharedReg333_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg333_out;
SharedReg899_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg899_out;
SharedReg105_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg105_out;
SharedReg726_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg726_out;
SharedReg1168_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1168_out;
SharedReg535_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg535_out;
SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg343_out;
SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg911_out;
SharedReg910_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg910_out;
SharedReg1429_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1429_out;
SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg345_out;
SharedReg334_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg334_out;
SharedReg901_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg901_out;
SharedReg99_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg99_out;
SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1155_out;
SharedReg913_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg913_out;
SharedReg87_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg87_out;
SharedReg713_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg713_out;
SharedReg543_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg543_out;
SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1155_out;
SharedReg349_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg349_out;
SharedReg95_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg95_out;
SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg921_out;
SharedReg355_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg355_out;
SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg921_out;
SharedReg1190_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1190_out;
SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg737_out;
SharedReg733_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg733_out;
SharedReg940_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg940_out;
SharedReg1191_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1191_out;
SharedReg548_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg548_out;
SharedReg124_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg124_out;
SharedReg950_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg950_out;
SharedReg382_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg382_out;
SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg737_out;
SharedReg1330_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1330_out;
SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg741_out;
SharedReg377_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg377_out;
SharedReg948_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg948_out;
SharedReg408_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg408_out;
SharedReg942_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg942_out;
   MUX_Subtract10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1354_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg552_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg3_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg17_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg6_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg11_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg16_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg333_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg899_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg105_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg726_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1168_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg535_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg97_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg911_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg910_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1429_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg345_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg334_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg901_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg99_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg913_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg87_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg713_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg543_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1155_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg349_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg95_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg355_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg921_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1190_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg569_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg733_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg940_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1191_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg548_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg124_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg950_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg382_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg737_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1330_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg741_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1196_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg377_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg948_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg408_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg942_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg549_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg348_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg100_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_3_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_0_out,
                 Y => Delay1No146_out);

SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg962_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg962_out;
SharedReg148_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg387_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
SharedReg1175_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1175_out;
SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg753_out;
SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg753_out;
SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg733_out;
SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg343_out;
SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg343_out;
SharedReg911_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg911_out;
SharedReg1430_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1430_out;
SharedReg1186_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1186_out;
SharedReg1181_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1181_out;
SharedReg1158_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1158_out;
SharedReg19_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg31_out;
SharedReg329_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg329_out;
SharedReg1360_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1360_out;
SharedReg107_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg107_out;
Delay41No20_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_27_cast <= Delay41No20_out;
SharedReg1171_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1171_out;
SharedReg725_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg725_out;
SharedReg109_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg109_out;
SharedReg924_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg924_out;
SharedReg938_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg938_out;
SharedReg1456_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1456_out;
SharedReg367_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg367_out;
SharedReg319_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg319_out;
SharedReg1431_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1431_out;
SharedReg338_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg338_out;
SharedReg1166_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1166_out;
SharedReg934_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg934_out;
SharedReg103_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg103_out;
SharedReg1160_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1160_out;
SharedReg1168_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1168_out;
SharedReg1161_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1161_out;
SharedReg344_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg344_out;
SharedReg349_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg349_out;
SharedReg910_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg910_out;
SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg95_out;
SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1428_out;
SharedReg747_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg747_out;
SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg733_out;
SharedReg1177_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1177_out;
SharedReg945_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg945_out;
SharedReg548_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg548_out;
SharedReg750_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg750_out;
SharedReg370_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg370_out;
SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1428_out;
SharedReg125_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg125_out;
SharedReg1193_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1193_out;
SharedReg949_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg949_out;
SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg748_out;
SharedReg153_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg153_out;
SharedReg1454_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1454_out;
SharedReg124_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg124_out;
SharedReg972_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg972_out;
   MUX_Subtract10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg962_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg911_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1430_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1186_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1181_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1158_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg19_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg21_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg35_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg24_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg148_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg34_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg31_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg329_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1360_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay41No20_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1171_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg725_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg109_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg387_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg924_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg938_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1456_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg367_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg319_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1431_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg338_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1166_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg934_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg103_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1175_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1160_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1168_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1161_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg344_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg349_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg910_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg95_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg747_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1177_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg945_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg548_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg750_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg370_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1428_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg125_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1193_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg949_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg753_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg153_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1454_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg124_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg972_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg733_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg343_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_3_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Subtract10_8_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Subtract10_8_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Subtract10_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_8_impl_out,
                 X => Delay1No148_out_to_Subtract10_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Subtract10_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg6_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg13_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg13_out;
SharedReg16_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg17_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg470_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg470_out;
SharedReg251_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg251_out;
SharedReg261_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg261_out;
SharedReg654_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg654_out;
SharedReg240_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg240_out;
SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg468_out;
SharedReg1104_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1104_out;
SharedReg467_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg467_out;
SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg657_out;
SharedReg1302_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1302_out;
SharedReg656_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg656_out;
SharedReg461_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg461_out;
SharedReg457_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg457_out;
SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1087_out;
SharedReg1093_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1093_out;
SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg657_out;
SharedReg477_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg477_out;
SharedReg1096_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1096_out;
SharedReg652_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg652_out;
SharedReg1474_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1474_out;
SharedReg473_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg473_out;
SharedReg1279_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1279_out;
SharedReg265_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_29_cast <= SharedReg265_out;
SharedReg661_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_30_cast <= SharedReg661_out;
SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_31_cast <= SharedReg841_out;
SharedReg465_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_32_cast <= SharedReg465_out;
SharedReg272_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_33_cast <= SharedReg272_out;
SharedReg837_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_34_cast <= SharedReg837_out;
SharedReg459_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_35_cast <= SharedReg459_out;
SharedReg1089_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1089_out;
SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1087_out;
SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1275_out;
SharedReg263_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_39_cast <= SharedReg263_out;
SharedReg1295_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1295_out;
SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1087_out;
SharedReg462_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_42_cast <= SharedReg462_out;
SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1275_out;
SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_44_cast <= SharedReg841_out;
SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1275_out;
SharedReg1464_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1464_out;
SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_47_cast <= SharedReg468_out;
SharedReg1097_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1097_out;
   MUX_Subtract10_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_48_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg240_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1104_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg467_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1302_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg656_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg461_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg457_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg6_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1093_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg657_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg477_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1096_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg652_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1474_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg473_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1279_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg265_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg661_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg13_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg465_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg272_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg837_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg459_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1089_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg263_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1295_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg16_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1087_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg462_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg841_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1275_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1464_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg468_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1097_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_48_cast,
                 iS_5 => SharedReg17_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg470_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg251_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg654_out_to_MUX_Subtract10_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract10_8_impl_0_LUT_out,
                 oMux => MUX_Subtract10_8_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_8_impl_0_out,
                 Y => Delay1No148_out);

SharedReg24_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg19_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg31_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg34_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg35_out;
SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg458_out;
SharedReg1095_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1095_out;
SharedReg235_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg235_out;
SharedReg1295_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1295_out;
SharedReg261_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg261_out;
SharedReg267_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg267_out;
SharedReg833_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg833_out;
SharedReg849_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg849_out;
SharedReg469_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg469_out;
SharedReg835_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg835_out;
SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg457_out;
SharedReg1087_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1087_out;
SharedReg262_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg262_out;
SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1281_out;
SharedReg1468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1468_out;
SharedReg243_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg243_out;
SharedReg1276_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1276_out;
SharedReg1089_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1089_out;
SharedReg1277_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1277_out;
SharedReg472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg472_out;
SharedReg468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg468_out;
SharedReg1086_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1086_out;
SharedReg1472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1472_out;
SharedReg1459_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1459_out;
SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_31_cast <= SharedReg457_out;
SharedReg1275_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1275_out;
SharedReg845_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_33_cast <= SharedReg845_out;
SharedReg286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_34_cast <= SharedReg286_out;
SharedReg289_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_35_cast <= SharedReg289_out;
SharedReg481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_36_cast <= SharedReg481_out;
SharedReg284_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_37_cast <= SharedReg284_out;
SharedReg1109_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1109_out;
SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1281_out;
SharedReg1293_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1293_out;
SharedReg1480_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1480_out;
SharedReg475_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_42_cast <= SharedReg475_out;
SharedReg1113_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1113_out;
SharedReg1278_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1278_out;
SharedReg1481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1481_out;
SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_46_cast <= SharedReg458_out;
SharedReg848_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_47_cast <= SharedReg848_out;
SharedReg1286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1286_out;
   MUX_Subtract10_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_48_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg261_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg267_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg833_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg849_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg469_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg835_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1087_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg262_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg243_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1276_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1089_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1277_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg468_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1086_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1472_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1459_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg31_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg457_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1275_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg845_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg289_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg284_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1109_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1281_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1293_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg34_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1480_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg475_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1113_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1278_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1481_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg848_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1286_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_48_cast,
                 iS_5 => SharedReg35_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg458_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1095_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1295_out_to_MUX_Subtract10_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract10_8_impl_1_LUT_out,
                 oMux => MUX_Subtract10_8_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_8_impl_1_out,
                 Y => Delay1No149_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay37No36_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => Delay37No36_out);

   Delay37No37_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => Delay37No37_out);

   Delay37No38_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => Delay37No38_out);

   Delay37No39_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => Delay37No39_out);

   Delay37No40_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => Delay37No40_out);

   Delay37No41_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => Delay37No41_out);

   Delay37No42_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => Delay37No42_out);

   Delay37No43_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => Delay37No43_out);

   Delay37No44_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => Delay37No44_out);

   Delay91No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay91No_out);

   Delay91No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay91No1_out);

   Delay91No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => Delay91No2_out);

   Delay91No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => Delay91No3_out);

   Delay91No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => Delay91No4_out);

   Delay91No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => Delay91No5_out);

   Delay91No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => Delay91No6_out);

   Delay91No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => Delay91No7_out);

   Delay91No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => Delay91No8_out);

   Delay43No9_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => Delay43No9_out);

   Delay43No10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => Delay43No10_out);

   Delay43No11_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => Delay43No11_out);

   Delay43No12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => Delay43No12_out);

   Delay43No13_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => Delay43No13_out);

   Delay43No14_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => Delay43No14_out);

   Delay43No15_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => Delay43No15_out);

   Delay43No16_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => Delay43No16_out);

   Delay43No17_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => Delay43No17_out);

   Delay41No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1134_out,
                 Y => Delay41No18_out);

   Delay41No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1154_out,
                 Y => Delay41No19_out);

   Delay41No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1174_out,
                 Y => Delay41No20_out);

   Delay41No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1194_out,
                 Y => Delay41No21_out);

   Delay41No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1214_out,
                 Y => Delay41No22_out);

   Delay41No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1234_out,
                 Y => Delay41No23_out);

   Delay41No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1254_out,
                 Y => Delay41No24_out);

   Delay41No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1274_out,
                 Y => Delay41No25_out);

   Delay41No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1294_out,
                 Y => Delay41No26_out);

   Delay80No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => Delay80No_out);

   Delay80No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => Delay80No1_out);

   Delay80No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => Delay80No2_out);

   Delay80No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => Delay80No3_out);

   Delay80No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => Delay80No4_out);

   Delay80No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => Delay80No6_out);

   Delay80No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => Delay80No8_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Add2_8_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add2_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_8_impl_0_LUT_out);

   MUX_Add2_8_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add2_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_8_impl_1_LUT_out);

   MUX_Add11_8_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add11_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add11_8_impl_0_LUT_out);

   MUX_Add11_8_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add11_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add11_8_impl_1_LUT_out);

   MUX_Subtract10_8_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract10_8_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract10_8_impl_0_LUT_out);

   MUX_Subtract10_8_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract10_8_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract10_8_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_5_impl_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_6_impl_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_7_impl_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_8_impl_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_5_impl_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_8_impl_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_5_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_6_impl_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_7_impl_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_8_impl_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_0_impl_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_1_impl_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_2_impl_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_3_impl_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_4_impl_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_5_impl_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_6_impl_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_7_impl_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_8_impl_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg857_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg918_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg934_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg938_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg965_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg971_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg983_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg984_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg985_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_5_impl_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1000_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1003_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1006_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1010_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);

   SharedReg1015_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => SharedReg1015_out);

   SharedReg1016_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1015_out,
                 Y => SharedReg1016_out);

   SharedReg1017_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1016_out,
                 Y => SharedReg1017_out);

   SharedReg1018_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1017_out,
                 Y => SharedReg1018_out);

   SharedReg1019_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1018_out,
                 Y => SharedReg1019_out);

   SharedReg1020_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1019_out,
                 Y => SharedReg1020_out);

   SharedReg1021_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1020_out,
                 Y => SharedReg1021_out);

   SharedReg1022_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1021_out,
                 Y => SharedReg1022_out);

   SharedReg1023_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1022_out,
                 Y => SharedReg1023_out);

   SharedReg1024_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1023_out,
                 Y => SharedReg1024_out);

   SharedReg1025_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1024_out,
                 Y => SharedReg1025_out);

   SharedReg1026_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1025_out,
                 Y => SharedReg1026_out);

   SharedReg1027_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_6_impl_out,
                 Y => SharedReg1027_out);

   SharedReg1028_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1027_out,
                 Y => SharedReg1028_out);

   SharedReg1029_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1028_out,
                 Y => SharedReg1029_out);

   SharedReg1030_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1029_out,
                 Y => SharedReg1030_out);

   SharedReg1031_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1030_out,
                 Y => SharedReg1031_out);

   SharedReg1032_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1031_out,
                 Y => SharedReg1032_out);

   SharedReg1033_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1032_out,
                 Y => SharedReg1033_out);

   SharedReg1034_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1033_out,
                 Y => SharedReg1034_out);

   SharedReg1035_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1034_out,
                 Y => SharedReg1035_out);

   SharedReg1036_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1035_out,
                 Y => SharedReg1036_out);

   SharedReg1037_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1036_out,
                 Y => SharedReg1037_out);

   SharedReg1038_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1037_out,
                 Y => SharedReg1038_out);

   SharedReg1039_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1038_out,
                 Y => SharedReg1039_out);

   SharedReg1040_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1039_out,
                 Y => SharedReg1040_out);

   SharedReg1041_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1040_out,
                 Y => SharedReg1041_out);

   SharedReg1042_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1041_out,
                 Y => SharedReg1042_out);

   SharedReg1043_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1042_out,
                 Y => SharedReg1043_out);

   SharedReg1044_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1043_out,
                 Y => SharedReg1044_out);

   SharedReg1045_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1044_out,
                 Y => SharedReg1045_out);

   SharedReg1046_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1045_out,
                 Y => SharedReg1046_out);

   SharedReg1047_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1046_out,
                 Y => SharedReg1047_out);

   SharedReg1048_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1047_out,
                 Y => SharedReg1048_out);

   SharedReg1049_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1048_out,
                 Y => SharedReg1049_out);

   SharedReg1050_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1049_out,
                 Y => SharedReg1050_out);

   SharedReg1051_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1050_out,
                 Y => SharedReg1051_out);

   SharedReg1052_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1051_out,
                 Y => SharedReg1052_out);

   SharedReg1053_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1052_out,
                 Y => SharedReg1053_out);

   SharedReg1054_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1053_out,
                 Y => SharedReg1054_out);

   SharedReg1055_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1054_out,
                 Y => SharedReg1055_out);

   SharedReg1056_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1055_out,
                 Y => SharedReg1056_out);

   SharedReg1057_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_7_impl_out,
                 Y => SharedReg1057_out);

   SharedReg1058_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1057_out,
                 Y => SharedReg1058_out);

   SharedReg1059_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1058_out,
                 Y => SharedReg1059_out);

   SharedReg1060_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1059_out,
                 Y => SharedReg1060_out);

   SharedReg1061_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1060_out,
                 Y => SharedReg1061_out);

   SharedReg1062_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1061_out,
                 Y => SharedReg1062_out);

   SharedReg1063_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1062_out,
                 Y => SharedReg1063_out);

   SharedReg1064_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1063_out,
                 Y => SharedReg1064_out);

   SharedReg1065_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1064_out,
                 Y => SharedReg1065_out);

   SharedReg1066_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1065_out,
                 Y => SharedReg1066_out);

   SharedReg1067_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1066_out,
                 Y => SharedReg1067_out);

   SharedReg1068_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1067_out,
                 Y => SharedReg1068_out);

   SharedReg1069_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1068_out,
                 Y => SharedReg1069_out);

   SharedReg1070_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1069_out,
                 Y => SharedReg1070_out);

   SharedReg1071_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1070_out,
                 Y => SharedReg1071_out);

   SharedReg1072_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1071_out,
                 Y => SharedReg1072_out);

   SharedReg1073_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1072_out,
                 Y => SharedReg1073_out);

   SharedReg1074_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1073_out,
                 Y => SharedReg1074_out);

   SharedReg1075_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1074_out,
                 Y => SharedReg1075_out);

   SharedReg1076_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1075_out,
                 Y => SharedReg1076_out);

   SharedReg1077_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1076_out,
                 Y => SharedReg1077_out);

   SharedReg1078_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1077_out,
                 Y => SharedReg1078_out);

   SharedReg1079_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1078_out,
                 Y => SharedReg1079_out);

   SharedReg1080_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1079_out,
                 Y => SharedReg1080_out);

   SharedReg1081_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1080_out,
                 Y => SharedReg1081_out);

   SharedReg1082_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1081_out,
                 Y => SharedReg1082_out);

   SharedReg1083_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1082_out,
                 Y => SharedReg1083_out);

   SharedReg1084_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1083_out,
                 Y => SharedReg1084_out);

   SharedReg1085_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1084_out,
                 Y => SharedReg1085_out);

   SharedReg1086_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_8_impl_out,
                 Y => SharedReg1086_out);

   SharedReg1087_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1086_out,
                 Y => SharedReg1087_out);

   SharedReg1088_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1087_out,
                 Y => SharedReg1088_out);

   SharedReg1089_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1088_out,
                 Y => SharedReg1089_out);

   SharedReg1090_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1089_out,
                 Y => SharedReg1090_out);

   SharedReg1091_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1090_out,
                 Y => SharedReg1091_out);

   SharedReg1092_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1091_out,
                 Y => SharedReg1092_out);

   SharedReg1093_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1092_out,
                 Y => SharedReg1093_out);

   SharedReg1094_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1093_out,
                 Y => SharedReg1094_out);

   SharedReg1095_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1094_out,
                 Y => SharedReg1095_out);

   SharedReg1096_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1095_out,
                 Y => SharedReg1096_out);

   SharedReg1097_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1096_out,
                 Y => SharedReg1097_out);

   SharedReg1098_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1097_out,
                 Y => SharedReg1098_out);

   SharedReg1099_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1098_out,
                 Y => SharedReg1099_out);

   SharedReg1100_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1099_out,
                 Y => SharedReg1100_out);

   SharedReg1101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1100_out,
                 Y => SharedReg1101_out);

   SharedReg1102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1101_out,
                 Y => SharedReg1102_out);

   SharedReg1103_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1102_out,
                 Y => SharedReg1103_out);

   SharedReg1104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1103_out,
                 Y => SharedReg1104_out);

   SharedReg1105_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1104_out,
                 Y => SharedReg1105_out);

   SharedReg1106_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1105_out,
                 Y => SharedReg1106_out);

   SharedReg1107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1106_out,
                 Y => SharedReg1107_out);

   SharedReg1108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1107_out,
                 Y => SharedReg1108_out);

   SharedReg1109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1108_out,
                 Y => SharedReg1109_out);

   SharedReg1110_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1109_out,
                 Y => SharedReg1110_out);

   SharedReg1111_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1110_out,
                 Y => SharedReg1111_out);

   SharedReg1112_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1111_out,
                 Y => SharedReg1112_out);

   SharedReg1113_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1112_out,
                 Y => SharedReg1113_out);

   SharedReg1114_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1113_out,
                 Y => SharedReg1114_out);

   SharedReg1115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg1115_out);

   SharedReg1116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1115_out,
                 Y => SharedReg1116_out);

   SharedReg1117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1116_out,
                 Y => SharedReg1117_out);

   SharedReg1118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1117_out,
                 Y => SharedReg1118_out);

   SharedReg1119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1118_out,
                 Y => SharedReg1119_out);

   SharedReg1120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1119_out,
                 Y => SharedReg1120_out);

   SharedReg1121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1120_out,
                 Y => SharedReg1121_out);

   SharedReg1122_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1121_out,
                 Y => SharedReg1122_out);

   SharedReg1123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1122_out,
                 Y => SharedReg1123_out);

   SharedReg1124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1123_out,
                 Y => SharedReg1124_out);

   SharedReg1125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1124_out,
                 Y => SharedReg1125_out);

   SharedReg1126_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1125_out,
                 Y => SharedReg1126_out);

   SharedReg1127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1126_out,
                 Y => SharedReg1127_out);

   SharedReg1128_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1127_out,
                 Y => SharedReg1128_out);

   SharedReg1129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1128_out,
                 Y => SharedReg1129_out);

   SharedReg1130_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1129_out,
                 Y => SharedReg1130_out);

   SharedReg1131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1130_out,
                 Y => SharedReg1131_out);

   SharedReg1132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1131_out,
                 Y => SharedReg1132_out);

   SharedReg1133_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1132_out,
                 Y => SharedReg1133_out);

   SharedReg1134_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1133_out,
                 Y => SharedReg1134_out);

   SharedReg1135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg1135_out);

   SharedReg1136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1135_out,
                 Y => SharedReg1136_out);

   SharedReg1137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1136_out,
                 Y => SharedReg1137_out);

   SharedReg1138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1137_out,
                 Y => SharedReg1138_out);

   SharedReg1139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1138_out,
                 Y => SharedReg1139_out);

   SharedReg1140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1139_out,
                 Y => SharedReg1140_out);

   SharedReg1141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1140_out,
                 Y => SharedReg1141_out);

   SharedReg1142_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1141_out,
                 Y => SharedReg1142_out);

   SharedReg1143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1142_out,
                 Y => SharedReg1143_out);

   SharedReg1144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1143_out,
                 Y => SharedReg1144_out);

   SharedReg1145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1144_out,
                 Y => SharedReg1145_out);

   SharedReg1146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1145_out,
                 Y => SharedReg1146_out);

   SharedReg1147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1146_out,
                 Y => SharedReg1147_out);

   SharedReg1148_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1147_out,
                 Y => SharedReg1148_out);

   SharedReg1149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1148_out,
                 Y => SharedReg1149_out);

   SharedReg1150_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1149_out,
                 Y => SharedReg1150_out);

   SharedReg1151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1150_out,
                 Y => SharedReg1151_out);

   SharedReg1152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1151_out,
                 Y => SharedReg1152_out);

   SharedReg1153_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1152_out,
                 Y => SharedReg1153_out);

   SharedReg1154_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1153_out,
                 Y => SharedReg1154_out);

   SharedReg1155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg1155_out);

   SharedReg1156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1155_out,
                 Y => SharedReg1156_out);

   SharedReg1157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1156_out,
                 Y => SharedReg1157_out);

   SharedReg1158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1157_out,
                 Y => SharedReg1158_out);

   SharedReg1159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1158_out,
                 Y => SharedReg1159_out);

   SharedReg1160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1159_out,
                 Y => SharedReg1160_out);

   SharedReg1161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1160_out,
                 Y => SharedReg1161_out);

   SharedReg1162_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1161_out,
                 Y => SharedReg1162_out);

   SharedReg1163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1162_out,
                 Y => SharedReg1163_out);

   SharedReg1164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1163_out,
                 Y => SharedReg1164_out);

   SharedReg1165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1164_out,
                 Y => SharedReg1165_out);

   SharedReg1166_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1165_out,
                 Y => SharedReg1166_out);

   SharedReg1167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1166_out,
                 Y => SharedReg1167_out);

   SharedReg1168_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1167_out,
                 Y => SharedReg1168_out);

   SharedReg1169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1168_out,
                 Y => SharedReg1169_out);

   SharedReg1170_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1169_out,
                 Y => SharedReg1170_out);

   SharedReg1171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1170_out,
                 Y => SharedReg1171_out);

   SharedReg1172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1171_out,
                 Y => SharedReg1172_out);

   SharedReg1173_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1172_out,
                 Y => SharedReg1173_out);

   SharedReg1174_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1173_out,
                 Y => SharedReg1174_out);

   SharedReg1175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg1175_out);

   SharedReg1176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1175_out,
                 Y => SharedReg1176_out);

   SharedReg1177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1176_out,
                 Y => SharedReg1177_out);

   SharedReg1178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1177_out,
                 Y => SharedReg1178_out);

   SharedReg1179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1178_out,
                 Y => SharedReg1179_out);

   SharedReg1180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1179_out,
                 Y => SharedReg1180_out);

   SharedReg1181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1180_out,
                 Y => SharedReg1181_out);

   SharedReg1182_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1181_out,
                 Y => SharedReg1182_out);

   SharedReg1183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1182_out,
                 Y => SharedReg1183_out);

   SharedReg1184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1183_out,
                 Y => SharedReg1184_out);

   SharedReg1185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1184_out,
                 Y => SharedReg1185_out);

   SharedReg1186_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1185_out,
                 Y => SharedReg1186_out);

   SharedReg1187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1186_out,
                 Y => SharedReg1187_out);

   SharedReg1188_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1187_out,
                 Y => SharedReg1188_out);

   SharedReg1189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1188_out,
                 Y => SharedReg1189_out);

   SharedReg1190_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1189_out,
                 Y => SharedReg1190_out);

   SharedReg1191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1190_out,
                 Y => SharedReg1191_out);

   SharedReg1192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1191_out,
                 Y => SharedReg1192_out);

   SharedReg1193_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1192_out,
                 Y => SharedReg1193_out);

   SharedReg1194_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1193_out,
                 Y => SharedReg1194_out);

   SharedReg1195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg1195_out);

   SharedReg1196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1195_out,
                 Y => SharedReg1196_out);

   SharedReg1197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1196_out,
                 Y => SharedReg1197_out);

   SharedReg1198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1197_out,
                 Y => SharedReg1198_out);

   SharedReg1199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1198_out,
                 Y => SharedReg1199_out);

   SharedReg1200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1199_out,
                 Y => SharedReg1200_out);

   SharedReg1201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1200_out,
                 Y => SharedReg1201_out);

   SharedReg1202_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1201_out,
                 Y => SharedReg1202_out);

   SharedReg1203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1202_out,
                 Y => SharedReg1203_out);

   SharedReg1204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1203_out,
                 Y => SharedReg1204_out);

   SharedReg1205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1204_out,
                 Y => SharedReg1205_out);

   SharedReg1206_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1205_out,
                 Y => SharedReg1206_out);

   SharedReg1207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1206_out,
                 Y => SharedReg1207_out);

   SharedReg1208_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1207_out,
                 Y => SharedReg1208_out);

   SharedReg1209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1208_out,
                 Y => SharedReg1209_out);

   SharedReg1210_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1209_out,
                 Y => SharedReg1210_out);

   SharedReg1211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1210_out,
                 Y => SharedReg1211_out);

   SharedReg1212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1211_out,
                 Y => SharedReg1212_out);

   SharedReg1213_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1212_out,
                 Y => SharedReg1213_out);

   SharedReg1214_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1213_out,
                 Y => SharedReg1214_out);

   SharedReg1215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_5_impl_out,
                 Y => SharedReg1215_out);

   SharedReg1216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1215_out,
                 Y => SharedReg1216_out);

   SharedReg1217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1216_out,
                 Y => SharedReg1217_out);

   SharedReg1218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1217_out,
                 Y => SharedReg1218_out);

   SharedReg1219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1218_out,
                 Y => SharedReg1219_out);

   SharedReg1220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1219_out,
                 Y => SharedReg1220_out);

   SharedReg1221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1220_out,
                 Y => SharedReg1221_out);

   SharedReg1222_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1221_out,
                 Y => SharedReg1222_out);

   SharedReg1223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1222_out,
                 Y => SharedReg1223_out);

   SharedReg1224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1223_out,
                 Y => SharedReg1224_out);

   SharedReg1225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1224_out,
                 Y => SharedReg1225_out);

   SharedReg1226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1225_out,
                 Y => SharedReg1226_out);

   SharedReg1227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1226_out,
                 Y => SharedReg1227_out);

   SharedReg1228_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1227_out,
                 Y => SharedReg1228_out);

   SharedReg1229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1228_out,
                 Y => SharedReg1229_out);

   SharedReg1230_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1229_out,
                 Y => SharedReg1230_out);

   SharedReg1231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1230_out,
                 Y => SharedReg1231_out);

   SharedReg1232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1231_out,
                 Y => SharedReg1232_out);

   SharedReg1233_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1232_out,
                 Y => SharedReg1233_out);

   SharedReg1234_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1233_out,
                 Y => SharedReg1234_out);

   SharedReg1235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_6_impl_out,
                 Y => SharedReg1235_out);

   SharedReg1236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1235_out,
                 Y => SharedReg1236_out);

   SharedReg1237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1236_out,
                 Y => SharedReg1237_out);

   SharedReg1238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1237_out,
                 Y => SharedReg1238_out);

   SharedReg1239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1238_out,
                 Y => SharedReg1239_out);

   SharedReg1240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1239_out,
                 Y => SharedReg1240_out);

   SharedReg1241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1240_out,
                 Y => SharedReg1241_out);

   SharedReg1242_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1241_out,
                 Y => SharedReg1242_out);

   SharedReg1243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1242_out,
                 Y => SharedReg1243_out);

   SharedReg1244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1243_out,
                 Y => SharedReg1244_out);

   SharedReg1245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1244_out,
                 Y => SharedReg1245_out);

   SharedReg1246_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1245_out,
                 Y => SharedReg1246_out);

   SharedReg1247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1246_out,
                 Y => SharedReg1247_out);

   SharedReg1248_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1247_out,
                 Y => SharedReg1248_out);

   SharedReg1249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1248_out,
                 Y => SharedReg1249_out);

   SharedReg1250_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1249_out,
                 Y => SharedReg1250_out);

   SharedReg1251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1250_out,
                 Y => SharedReg1251_out);

   SharedReg1252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1251_out,
                 Y => SharedReg1252_out);

   SharedReg1253_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1252_out,
                 Y => SharedReg1253_out);

   SharedReg1254_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1253_out,
                 Y => SharedReg1254_out);

   SharedReg1255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_7_impl_out,
                 Y => SharedReg1255_out);

   SharedReg1256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1255_out,
                 Y => SharedReg1256_out);

   SharedReg1257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1256_out,
                 Y => SharedReg1257_out);

   SharedReg1258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1257_out,
                 Y => SharedReg1258_out);

   SharedReg1259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1258_out,
                 Y => SharedReg1259_out);

   SharedReg1260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1259_out,
                 Y => SharedReg1260_out);

   SharedReg1261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1260_out,
                 Y => SharedReg1261_out);

   SharedReg1262_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1261_out,
                 Y => SharedReg1262_out);

   SharedReg1263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1262_out,
                 Y => SharedReg1263_out);

   SharedReg1264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1263_out,
                 Y => SharedReg1264_out);

   SharedReg1265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1264_out,
                 Y => SharedReg1265_out);

   SharedReg1266_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1265_out,
                 Y => SharedReg1266_out);

   SharedReg1267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1266_out,
                 Y => SharedReg1267_out);

   SharedReg1268_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1267_out,
                 Y => SharedReg1268_out);

   SharedReg1269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1268_out,
                 Y => SharedReg1269_out);

   SharedReg1270_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1269_out,
                 Y => SharedReg1270_out);

   SharedReg1271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1270_out,
                 Y => SharedReg1271_out);

   SharedReg1272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1271_out,
                 Y => SharedReg1272_out);

   SharedReg1273_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1272_out,
                 Y => SharedReg1273_out);

   SharedReg1274_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1273_out,
                 Y => SharedReg1274_out);

   SharedReg1275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_8_impl_out,
                 Y => SharedReg1275_out);

   SharedReg1276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1275_out,
                 Y => SharedReg1276_out);

   SharedReg1277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1276_out,
                 Y => SharedReg1277_out);

   SharedReg1278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1277_out,
                 Y => SharedReg1278_out);

   SharedReg1279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1278_out,
                 Y => SharedReg1279_out);

   SharedReg1280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1279_out,
                 Y => SharedReg1280_out);

   SharedReg1281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1280_out,
                 Y => SharedReg1281_out);

   SharedReg1282_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1281_out,
                 Y => SharedReg1282_out);

   SharedReg1283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1282_out,
                 Y => SharedReg1283_out);

   SharedReg1284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1283_out,
                 Y => SharedReg1284_out);

   SharedReg1285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1284_out,
                 Y => SharedReg1285_out);

   SharedReg1286_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1285_out,
                 Y => SharedReg1286_out);

   SharedReg1287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1286_out,
                 Y => SharedReg1287_out);

   SharedReg1288_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1287_out,
                 Y => SharedReg1288_out);

   SharedReg1289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1288_out,
                 Y => SharedReg1289_out);

   SharedReg1290_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1289_out,
                 Y => SharedReg1290_out);

   SharedReg1291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1290_out,
                 Y => SharedReg1291_out);

   SharedReg1292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1291_out,
                 Y => SharedReg1292_out);

   SharedReg1293_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1292_out,
                 Y => SharedReg1293_out);

   SharedReg1294_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1293_out,
                 Y => SharedReg1294_out);

   SharedReg1295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_8_impl_out,
                 Y => SharedReg1295_out);

   SharedReg1296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1295_out,
                 Y => SharedReg1296_out);

   SharedReg1297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1296_out,
                 Y => SharedReg1297_out);

   SharedReg1298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1297_out,
                 Y => SharedReg1298_out);

   SharedReg1299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1298_out,
                 Y => SharedReg1299_out);

   SharedReg1300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1299_out,
                 Y => SharedReg1300_out);

   SharedReg1301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1300_out,
                 Y => SharedReg1301_out);

   SharedReg1302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1301_out,
                 Y => SharedReg1302_out);

   SharedReg1303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1302_out,
                 Y => SharedReg1303_out);

   SharedReg1304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1303_out,
                 Y => SharedReg1304_out);

   SharedReg1305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1304_out,
                 Y => SharedReg1305_out);

   SharedReg1306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1305_out,
                 Y => SharedReg1306_out);

   SharedReg1307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1306_out,
                 Y => SharedReg1307_out);

   SharedReg1308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1307_out,
                 Y => SharedReg1308_out);

   SharedReg1309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1308_out,
                 Y => SharedReg1309_out);

   SharedReg1310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1309_out,
                 Y => SharedReg1310_out);

   SharedReg1311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1310_out,
                 Y => SharedReg1311_out);

   SharedReg1312_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1311_out,
                 Y => SharedReg1312_out);

   SharedReg1313_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1312_out,
                 Y => SharedReg1313_out);

   SharedReg1314_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1313_out,
                 Y => SharedReg1314_out);

   SharedReg1315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1314_out,
                 Y => SharedReg1315_out);

   SharedReg1316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1315_out,
                 Y => SharedReg1316_out);

   SharedReg1317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1316_out,
                 Y => SharedReg1317_out);

   SharedReg1318_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1317_out,
                 Y => SharedReg1318_out);

   SharedReg1319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1318_out,
                 Y => SharedReg1319_out);

   SharedReg1320_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1319_out,
                 Y => SharedReg1320_out);

   SharedReg1321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_4_impl_out,
                 Y => SharedReg1321_out);

   SharedReg1322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1321_out,
                 Y => SharedReg1322_out);

   SharedReg1323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1322_out,
                 Y => SharedReg1323_out);

   SharedReg1324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1323_out,
                 Y => SharedReg1324_out);

   SharedReg1325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1324_out,
                 Y => SharedReg1325_out);

   SharedReg1326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1325_out,
                 Y => SharedReg1326_out);

   SharedReg1327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1326_out,
                 Y => SharedReg1327_out);

   SharedReg1328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1327_out,
                 Y => SharedReg1328_out);

   SharedReg1329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1328_out,
                 Y => SharedReg1329_out);

   SharedReg1330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1329_out,
                 Y => SharedReg1330_out);

   SharedReg1331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1330_out,
                 Y => SharedReg1331_out);

   SharedReg1332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1331_out,
                 Y => SharedReg1332_out);

   SharedReg1333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1332_out,
                 Y => SharedReg1333_out);

   SharedReg1334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1333_out,
                 Y => SharedReg1334_out);

   SharedReg1335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1334_out,
                 Y => SharedReg1335_out);

   SharedReg1336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1335_out,
                 Y => SharedReg1336_out);

   SharedReg1337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1336_out,
                 Y => SharedReg1337_out);

   SharedReg1338_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1337_out,
                 Y => SharedReg1338_out);

   SharedReg1339_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1338_out,
                 Y => SharedReg1339_out);

   SharedReg1340_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1339_out,
                 Y => SharedReg1340_out);

   SharedReg1341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1340_out,
                 Y => SharedReg1341_out);

   SharedReg1342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1341_out,
                 Y => SharedReg1342_out);

   SharedReg1343_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1342_out,
                 Y => SharedReg1343_out);

   SharedReg1344_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1343_out,
                 Y => SharedReg1344_out);

   SharedReg1345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1344_out,
                 Y => SharedReg1345_out);

   SharedReg1346_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1345_out,
                 Y => SharedReg1346_out);

   SharedReg1347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_2_impl_out,
                 Y => SharedReg1347_out);

   SharedReg1348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1347_out,
                 Y => SharedReg1348_out);

   SharedReg1349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1348_out,
                 Y => SharedReg1349_out);

   SharedReg1350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1349_out,
                 Y => SharedReg1350_out);

   SharedReg1351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1350_out,
                 Y => SharedReg1351_out);

   SharedReg1352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1351_out,
                 Y => SharedReg1352_out);

   SharedReg1353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1352_out,
                 Y => SharedReg1353_out);

   SharedReg1354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1353_out,
                 Y => SharedReg1354_out);

   SharedReg1355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1354_out,
                 Y => SharedReg1355_out);

   SharedReg1356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1355_out,
                 Y => SharedReg1356_out);

   SharedReg1357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1356_out,
                 Y => SharedReg1357_out);

   SharedReg1358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1357_out,
                 Y => SharedReg1358_out);

   SharedReg1359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1358_out,
                 Y => SharedReg1359_out);

   SharedReg1360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1359_out,
                 Y => SharedReg1360_out);

   SharedReg1361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1360_out,
                 Y => SharedReg1361_out);

   SharedReg1362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1361_out,
                 Y => SharedReg1362_out);

   SharedReg1363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1362_out,
                 Y => SharedReg1363_out);

   SharedReg1364_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1363_out,
                 Y => SharedReg1364_out);

   SharedReg1365_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1364_out,
                 Y => SharedReg1365_out);

   SharedReg1366_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1365_out,
                 Y => SharedReg1366_out);

   SharedReg1367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1366_out,
                 Y => SharedReg1367_out);

   SharedReg1368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1367_out,
                 Y => SharedReg1368_out);

   SharedReg1369_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1368_out,
                 Y => SharedReg1369_out);

   SharedReg1370_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1369_out,
                 Y => SharedReg1370_out);

   SharedReg1371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1370_out,
                 Y => SharedReg1371_out);

   SharedReg1372_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1371_out,
                 Y => SharedReg1372_out);

   SharedReg1373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_7_impl_out,
                 Y => SharedReg1373_out);

   SharedReg1374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1373_out,
                 Y => SharedReg1374_out);

   SharedReg1375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1374_out,
                 Y => SharedReg1375_out);

   SharedReg1376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1375_out,
                 Y => SharedReg1376_out);

   SharedReg1377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1376_out,
                 Y => SharedReg1377_out);

   SharedReg1378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1377_out,
                 Y => SharedReg1378_out);

   SharedReg1379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1378_out,
                 Y => SharedReg1379_out);

   SharedReg1380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1379_out,
                 Y => SharedReg1380_out);

   SharedReg1381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1380_out,
                 Y => SharedReg1381_out);

   SharedReg1382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1381_out,
                 Y => SharedReg1382_out);

   SharedReg1383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1382_out,
                 Y => SharedReg1383_out);

   SharedReg1384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1383_out,
                 Y => SharedReg1384_out);

   SharedReg1385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1384_out,
                 Y => SharedReg1385_out);

   SharedReg1386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1385_out,
                 Y => SharedReg1386_out);

   SharedReg1387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1386_out,
                 Y => SharedReg1387_out);

   SharedReg1388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1387_out,
                 Y => SharedReg1388_out);

   SharedReg1389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1388_out,
                 Y => SharedReg1389_out);

   SharedReg1390_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1389_out,
                 Y => SharedReg1390_out);

   SharedReg1391_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1390_out,
                 Y => SharedReg1391_out);

   SharedReg1392_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1391_out,
                 Y => SharedReg1392_out);

   SharedReg1393_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1392_out,
                 Y => SharedReg1393_out);

   SharedReg1394_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1393_out,
                 Y => SharedReg1394_out);

   SharedReg1395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1394_out,
                 Y => SharedReg1395_out);

   SharedReg1396_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1395_out,
                 Y => SharedReg1396_out);

   SharedReg1397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1396_out,
                 Y => SharedReg1397_out);

   SharedReg1398_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1397_out,
                 Y => SharedReg1398_out);

   SharedReg1399_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1398_out,
                 Y => SharedReg1399_out);

   SharedReg1400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_1_impl_out,
                 Y => SharedReg1400_out);

   SharedReg1401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1400_out,
                 Y => SharedReg1401_out);

   SharedReg1402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1401_out,
                 Y => SharedReg1402_out);

   SharedReg1403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1402_out,
                 Y => SharedReg1403_out);

   SharedReg1404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1403_out,
                 Y => SharedReg1404_out);

   SharedReg1405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1404_out,
                 Y => SharedReg1405_out);

   SharedReg1406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1405_out,
                 Y => SharedReg1406_out);

   SharedReg1407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1406_out,
                 Y => SharedReg1407_out);

   SharedReg1408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1407_out,
                 Y => SharedReg1408_out);

   SharedReg1409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1408_out,
                 Y => SharedReg1409_out);

   SharedReg1410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1409_out,
                 Y => SharedReg1410_out);

   SharedReg1411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1410_out,
                 Y => SharedReg1411_out);

   SharedReg1412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1411_out,
                 Y => SharedReg1412_out);

   SharedReg1413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1412_out,
                 Y => SharedReg1413_out);

   SharedReg1414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1413_out,
                 Y => SharedReg1414_out);

   SharedReg1415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1414_out,
                 Y => SharedReg1415_out);

   SharedReg1416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1415_out,
                 Y => SharedReg1416_out);

   SharedReg1417_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1416_out,
                 Y => SharedReg1417_out);

   SharedReg1418_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1417_out,
                 Y => SharedReg1418_out);

   SharedReg1419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1418_out,
                 Y => SharedReg1419_out);

   SharedReg1420_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1419_out,
                 Y => SharedReg1420_out);

   SharedReg1421_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1420_out,
                 Y => SharedReg1421_out);

   SharedReg1422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1421_out,
                 Y => SharedReg1422_out);

   SharedReg1423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1422_out,
                 Y => SharedReg1423_out);

   SharedReg1424_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1423_out,
                 Y => SharedReg1424_out);

   SharedReg1425_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1424_out,
                 Y => SharedReg1425_out);

   SharedReg1426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1425_out,
                 Y => SharedReg1426_out);

   SharedReg1427_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1426_out,
                 Y => SharedReg1427_out);

   SharedReg1428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_3_impl_out,
                 Y => SharedReg1428_out);

   SharedReg1429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1428_out,
                 Y => SharedReg1429_out);

   SharedReg1430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1429_out,
                 Y => SharedReg1430_out);

   SharedReg1431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1430_out,
                 Y => SharedReg1431_out);

   SharedReg1432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1431_out,
                 Y => SharedReg1432_out);

   SharedReg1433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1432_out,
                 Y => SharedReg1433_out);

   SharedReg1434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1433_out,
                 Y => SharedReg1434_out);

   SharedReg1435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1434_out,
                 Y => SharedReg1435_out);

   SharedReg1436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1435_out,
                 Y => SharedReg1436_out);

   SharedReg1437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1436_out,
                 Y => SharedReg1437_out);

   SharedReg1438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1437_out,
                 Y => SharedReg1438_out);

   SharedReg1439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1438_out,
                 Y => SharedReg1439_out);

   SharedReg1440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1439_out,
                 Y => SharedReg1440_out);

   SharedReg1441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1440_out,
                 Y => SharedReg1441_out);

   SharedReg1442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1441_out,
                 Y => SharedReg1442_out);

   SharedReg1443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1442_out,
                 Y => SharedReg1443_out);

   SharedReg1444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1443_out,
                 Y => SharedReg1444_out);

   SharedReg1445_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1444_out,
                 Y => SharedReg1445_out);

   SharedReg1446_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1445_out,
                 Y => SharedReg1446_out);

   SharedReg1447_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1446_out,
                 Y => SharedReg1447_out);

   SharedReg1448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1447_out,
                 Y => SharedReg1448_out);

   SharedReg1449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1448_out,
                 Y => SharedReg1449_out);

   SharedReg1450_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1449_out,
                 Y => SharedReg1450_out);

   SharedReg1451_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1450_out,
                 Y => SharedReg1451_out);

   SharedReg1452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1451_out,
                 Y => SharedReg1452_out);

   SharedReg1453_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1452_out,
                 Y => SharedReg1453_out);

   SharedReg1454_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1453_out,
                 Y => SharedReg1454_out);

   SharedReg1455_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1454_out,
                 Y => SharedReg1455_out);

   SharedReg1456_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1455_out,
                 Y => SharedReg1456_out);

   SharedReg1457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_8_impl_out,
                 Y => SharedReg1457_out);

   SharedReg1458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1457_out,
                 Y => SharedReg1458_out);

   SharedReg1459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1458_out,
                 Y => SharedReg1459_out);

   SharedReg1460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1459_out,
                 Y => SharedReg1460_out);

   SharedReg1461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1460_out,
                 Y => SharedReg1461_out);

   SharedReg1462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1461_out,
                 Y => SharedReg1462_out);

   SharedReg1463_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1462_out,
                 Y => SharedReg1463_out);

   SharedReg1464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1463_out,
                 Y => SharedReg1464_out);

   SharedReg1465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1464_out,
                 Y => SharedReg1465_out);

   SharedReg1466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1465_out,
                 Y => SharedReg1466_out);

   SharedReg1467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1466_out,
                 Y => SharedReg1467_out);

   SharedReg1468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1467_out,
                 Y => SharedReg1468_out);

   SharedReg1469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1468_out,
                 Y => SharedReg1469_out);

   SharedReg1470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1469_out,
                 Y => SharedReg1470_out);

   SharedReg1471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1470_out,
                 Y => SharedReg1471_out);

   SharedReg1472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1471_out,
                 Y => SharedReg1472_out);

   SharedReg1473_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1472_out,
                 Y => SharedReg1473_out);

   SharedReg1474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1473_out,
                 Y => SharedReg1474_out);

   SharedReg1475_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1474_out,
                 Y => SharedReg1475_out);

   SharedReg1476_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1475_out,
                 Y => SharedReg1476_out);

   SharedReg1477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1476_out,
                 Y => SharedReg1477_out);

   SharedReg1478_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1477_out,
                 Y => SharedReg1478_out);

   SharedReg1479_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1478_out,
                 Y => SharedReg1479_out);

   SharedReg1480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1479_out,
                 Y => SharedReg1480_out);

   SharedReg1481_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1480_out,
                 Y => SharedReg1481_out);

   SharedReg1482_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg1482_out);

   SharedReg1483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1482_out,
                 Y => SharedReg1483_out);

   SharedReg1484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1483_out,
                 Y => SharedReg1484_out);

   SharedReg1485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1484_out,
                 Y => SharedReg1485_out);

   SharedReg1486_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1485_out,
                 Y => SharedReg1486_out);

   SharedReg1487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1486_out,
                 Y => SharedReg1487_out);

   SharedReg1488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1487_out,
                 Y => SharedReg1488_out);

   SharedReg1489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1488_out,
                 Y => SharedReg1489_out);

   SharedReg1490_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1489_out,
                 Y => SharedReg1490_out);

   SharedReg1491_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1490_out,
                 Y => SharedReg1491_out);

   SharedReg1492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1491_out,
                 Y => SharedReg1492_out);

   SharedReg1493_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1492_out,
                 Y => SharedReg1493_out);

   SharedReg1494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1493_out,
                 Y => SharedReg1494_out);

   SharedReg1495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1494_out,
                 Y => SharedReg1495_out);

   SharedReg1496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1495_out,
                 Y => SharedReg1496_out);

   SharedReg1497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1496_out,
                 Y => SharedReg1497_out);

   SharedReg1498_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1497_out,
                 Y => SharedReg1498_out);

   SharedReg1499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1498_out,
                 Y => SharedReg1499_out);

   SharedReg1500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1499_out,
                 Y => SharedReg1500_out);

   SharedReg1501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1500_out,
                 Y => SharedReg1501_out);

   SharedReg1502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1501_out,
                 Y => SharedReg1502_out);

   SharedReg1503_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1502_out,
                 Y => SharedReg1503_out);

   SharedReg1504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1503_out,
                 Y => SharedReg1504_out);

   SharedReg1505_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1504_out,
                 Y => SharedReg1505_out);

   SharedReg1506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1505_out,
                 Y => SharedReg1506_out);

   SharedReg1507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1506_out,
                 Y => SharedReg1507_out);

   SharedReg1508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1507_out,
                 Y => SharedReg1508_out);

   SharedReg1509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1508_out,
                 Y => SharedReg1509_out);

   SharedReg1510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1509_out,
                 Y => SharedReg1510_out);

   SharedReg1511_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1510_out,
                 Y => SharedReg1511_out);

   SharedReg1512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1511_out,
                 Y => SharedReg1512_out);

   SharedReg1513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1512_out,
                 Y => SharedReg1513_out);

   SharedReg1514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1513_out,
                 Y => SharedReg1514_out);

   SharedReg1515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1514_out,
                 Y => SharedReg1515_out);

   SharedReg1516_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1515_out,
                 Y => SharedReg1516_out);

   SharedReg1517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1516_out,
                 Y => SharedReg1517_out);

   SharedReg1518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1517_out,
                 Y => SharedReg1518_out);

   SharedReg1519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1518_out,
                 Y => SharedReg1519_out);

   SharedReg1520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1519_out,
                 Y => SharedReg1520_out);

   SharedReg1521_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1520_out,
                 Y => SharedReg1521_out);

   SharedReg1522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1521_out,
                 Y => SharedReg1522_out);

   SharedReg1523_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1522_out,
                 Y => SharedReg1523_out);

   SharedReg1524_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1523_out,
                 Y => SharedReg1524_out);

   SharedReg1525_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1524_out,
                 Y => SharedReg1525_out);

   SharedReg1526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1525_out,
                 Y => SharedReg1526_out);

   SharedReg1527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1526_out,
                 Y => SharedReg1527_out);

   SharedReg1528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1527_out,
                 Y => SharedReg1528_out);

   SharedReg1529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1528_out,
                 Y => SharedReg1529_out);

   SharedReg1530_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1529_out,
                 Y => SharedReg1530_out);

   SharedReg1531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1530_out,
                 Y => SharedReg1531_out);

   SharedReg1532_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1531_out,
                 Y => SharedReg1532_out);

   SharedReg1533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1532_out,
                 Y => SharedReg1533_out);

   SharedReg1534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1533_out,
                 Y => SharedReg1534_out);

   SharedReg1535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1534_out,
                 Y => SharedReg1535_out);

   SharedReg1536_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1535_out,
                 Y => SharedReg1536_out);

   SharedReg1537_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg1537_out);

   SharedReg1538_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1537_out,
                 Y => SharedReg1538_out);

   SharedReg1539_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1538_out,
                 Y => SharedReg1539_out);

   SharedReg1540_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1539_out,
                 Y => SharedReg1540_out);

   SharedReg1541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1540_out,
                 Y => SharedReg1541_out);

   SharedReg1542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1541_out,
                 Y => SharedReg1542_out);

   SharedReg1543_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1542_out,
                 Y => SharedReg1543_out);

   SharedReg1544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1543_out,
                 Y => SharedReg1544_out);

   SharedReg1545_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1544_out,
                 Y => SharedReg1545_out);

   SharedReg1546_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1545_out,
                 Y => SharedReg1546_out);

   SharedReg1547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1546_out,
                 Y => SharedReg1547_out);

   SharedReg1548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1547_out,
                 Y => SharedReg1548_out);

   SharedReg1549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1548_out,
                 Y => SharedReg1549_out);

   SharedReg1550_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1549_out,
                 Y => SharedReg1550_out);

   SharedReg1551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1550_out,
                 Y => SharedReg1551_out);

   SharedReg1552_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1551_out,
                 Y => SharedReg1552_out);

   SharedReg1553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1552_out,
                 Y => SharedReg1553_out);

   SharedReg1554_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1553_out,
                 Y => SharedReg1554_out);

   SharedReg1555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1554_out,
                 Y => SharedReg1555_out);

   SharedReg1556_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1555_out,
                 Y => SharedReg1556_out);

   SharedReg1557_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1556_out,
                 Y => SharedReg1557_out);

   SharedReg1558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1557_out,
                 Y => SharedReg1558_out);

   SharedReg1559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1558_out,
                 Y => SharedReg1559_out);

   SharedReg1560_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1559_out,
                 Y => SharedReg1560_out);

   SharedReg1561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1560_out,
                 Y => SharedReg1561_out);

   SharedReg1562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1561_out,
                 Y => SharedReg1562_out);

   SharedReg1563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1562_out,
                 Y => SharedReg1563_out);

   SharedReg1564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1563_out,
                 Y => SharedReg1564_out);

   SharedReg1565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1564_out,
                 Y => SharedReg1565_out);

   SharedReg1566_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1565_out,
                 Y => SharedReg1566_out);

   SharedReg1567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1566_out,
                 Y => SharedReg1567_out);

   SharedReg1568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1567_out,
                 Y => SharedReg1568_out);

   SharedReg1569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1568_out,
                 Y => SharedReg1569_out);

   SharedReg1570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1569_out,
                 Y => SharedReg1570_out);

   SharedReg1571_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1570_out,
                 Y => SharedReg1571_out);

   SharedReg1572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1571_out,
                 Y => SharedReg1572_out);

   SharedReg1573_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1572_out,
                 Y => SharedReg1573_out);

   SharedReg1574_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1573_out,
                 Y => SharedReg1574_out);

   SharedReg1575_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1574_out,
                 Y => SharedReg1575_out);

   SharedReg1576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1575_out,
                 Y => SharedReg1576_out);

   SharedReg1577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1576_out,
                 Y => SharedReg1577_out);

   SharedReg1578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1577_out,
                 Y => SharedReg1578_out);

   SharedReg1579_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1578_out,
                 Y => SharedReg1579_out);

   SharedReg1580_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1579_out,
                 Y => SharedReg1580_out);

   SharedReg1581_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1580_out,
                 Y => SharedReg1581_out);

   SharedReg1582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1581_out,
                 Y => SharedReg1582_out);

   SharedReg1583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1582_out,
                 Y => SharedReg1583_out);

   SharedReg1584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1583_out,
                 Y => SharedReg1584_out);

   SharedReg1585_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1584_out,
                 Y => SharedReg1585_out);

   SharedReg1586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1585_out,
                 Y => SharedReg1586_out);

   SharedReg1587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1586_out,
                 Y => SharedReg1587_out);

   SharedReg1588_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg1588_out);

   SharedReg1589_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1588_out,
                 Y => SharedReg1589_out);

   SharedReg1590_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1589_out,
                 Y => SharedReg1590_out);

   SharedReg1591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1590_out,
                 Y => SharedReg1591_out);

   SharedReg1592_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1591_out,
                 Y => SharedReg1592_out);

   SharedReg1593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1592_out,
                 Y => SharedReg1593_out);

   SharedReg1594_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg1594_out);

   SharedReg1595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1594_out,
                 Y => SharedReg1595_out);

   SharedReg1596_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1595_out,
                 Y => SharedReg1596_out);

   SharedReg1597_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1596_out,
                 Y => SharedReg1597_out);

   SharedReg1598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1597_out,
                 Y => SharedReg1598_out);

   SharedReg1599_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1598_out,
                 Y => SharedReg1599_out);

   SharedReg1600_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg1600_out);

   SharedReg1601_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg1601_out);

   SharedReg1602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1601_out,
                 Y => SharedReg1602_out);

   SharedReg1603_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg1603_out);

   SharedReg1604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1603_out,
                 Y => SharedReg1604_out);

   SharedReg1605_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1604_out,
                 Y => SharedReg1605_out);

   SharedReg1606_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1605_out,
                 Y => SharedReg1606_out);

   SharedReg1607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1606_out,
                 Y => SharedReg1607_out);

   SharedReg1608_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1607_out,
                 Y => SharedReg1608_out);

   SharedReg1609_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1608_out,
                 Y => SharedReg1609_out);

   SharedReg1610_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1609_out,
                 Y => SharedReg1610_out);

   SharedReg1611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1610_out,
                 Y => SharedReg1611_out);

   SharedReg1612_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1611_out,
                 Y => SharedReg1612_out);

   SharedReg1613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1612_out,
                 Y => SharedReg1613_out);

   SharedReg1614_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1613_out,
                 Y => SharedReg1614_out);

   SharedReg1615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1614_out,
                 Y => SharedReg1615_out);

   SharedReg1616_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg1616_out);

   SharedReg1617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1616_out,
                 Y => SharedReg1617_out);

   SharedReg1618_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1617_out,
                 Y => SharedReg1618_out);

   SharedReg1619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1618_out,
                 Y => SharedReg1619_out);

   SharedReg1620_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1619_out,
                 Y => SharedReg1620_out);

   SharedReg1621_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1620_out,
                 Y => SharedReg1621_out);

   SharedReg1622_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1621_out,
                 Y => SharedReg1622_out);

   SharedReg1623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1622_out,
                 Y => SharedReg1623_out);

   SharedReg1624_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1623_out,
                 Y => SharedReg1624_out);

   SharedReg1625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1624_out,
                 Y => SharedReg1625_out);

   SharedReg1626_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1625_out,
                 Y => SharedReg1626_out);

   SharedReg1627_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1626_out,
                 Y => SharedReg1627_out);

   SharedReg1628_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1627_out,
                 Y => SharedReg1628_out);

   SharedReg1629_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1628_out,
                 Y => SharedReg1629_out);

   SharedReg1630_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg1630_out);

   SharedReg1631_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1630_out,
                 Y => SharedReg1631_out);

   SharedReg1632_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg1632_out);

   SharedReg1633_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1632_out,
                 Y => SharedReg1633_out);

   SharedReg1634_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg1634_out);

   SharedReg1635_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1634_out,
                 Y => SharedReg1635_out);

   SharedReg1636_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1635_out,
                 Y => SharedReg1636_out);

   SharedReg1637_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1636_out,
                 Y => SharedReg1637_out);

   SharedReg1638_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1637_out,
                 Y => SharedReg1638_out);

   SharedReg1639_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1638_out,
                 Y => SharedReg1639_out);

   SharedReg1640_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg1640_out);

   SharedReg1641_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1640_out,
                 Y => SharedReg1641_out);

   SharedReg1642_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1641_out,
                 Y => SharedReg1642_out);

   SharedReg1643_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1642_out,
                 Y => SharedReg1643_out);

   SharedReg1644_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1643_out,
                 Y => SharedReg1644_out);

   SharedReg1645_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1644_out,
                 Y => SharedReg1645_out);

   SharedReg1646_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg1646_out);

   SharedReg1647_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1646_out,
                 Y => SharedReg1647_out);

   SharedReg1648_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg1648_out);

   SharedReg1649_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1648_out,
                 Y => SharedReg1649_out);

   SharedReg1650_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg1650_out);

   SharedReg1651_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg1651_out);
end architecture;

