--------------------------------------------------------------------------------
--                         ModuloCounter_14_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_14_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_14_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 13 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1668762
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1668762 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1668762 is
signal XX_m1668763 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1668763 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1668763 <= X ;
   YY_m1668763 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1668766
--                   (IntAdderClassical_33_f500_uid1668768)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1668766 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1668766 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1668762 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1668766 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1668762  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid1668766  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_14_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_14_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_14_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
         iS_13 when "1101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1669757_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1669759)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1669757_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1669757_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1669762
--                  (IntAdderAlternative_27_f250_uid1669766)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1669762 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1669762 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1669769
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1669769 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1669769 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1669772
--                   (IntAdderClassical_34_f250_uid1669774)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1669772 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1669772 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1669757
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1669757 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1669757 is
   component FPAdd_8_23_uid1669757_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1669762 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1669769 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1669772 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1669757_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1669762  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1669769  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1669772  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1669757 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1669757  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_7_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_12_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1670813_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1670815)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1670813_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1670813_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1670818
--                  (IntAdderAlternative_27_f250_uid1670822)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1670818 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1670818 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1670825
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1670825 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1670825 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1670828
--                   (IntAdderClassical_34_f250_uid1670830)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1670828 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1670828 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1670813
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1670813 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1670813 is
   component FPAdd_8_23_uid1670813_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1670818 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1670825 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1670828 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1670813_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1670818  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1670825  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1670828  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid1670813 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid1670813  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_9_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_133_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 133 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_133_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_133_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      Y <= s132;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 139 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      Y <= s138;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      Y <= s40;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      Y <= s62;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      Y <= s55;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 80 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      Y <= s79;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 122 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      Y <= s121;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 96 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      Y <= s95;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 40 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      Y <= s39;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 115 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      Y <= s114;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 45 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      Y <= s44;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "010" when "0000",
      "110" when "0001",
      "000" when "0010",
      "011" when "0011",
      "000" when "0100",
      "000" when "0101",
      "101" when "0110",
      "000" when "0111",
      "000" when "1000",
      "001" when "1001",
      "000" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "010" when "0000",
      "011" when "0001",
      "000" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "000" when "1000",
      "000" when "1001",
      "000" when "1010",
      "001" when "1011",
      "101" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "1011" when "0000",
      "0101" when "0001",
      "1001" when "0010",
      "0111" when "0011",
      "0011" when "0100",
      "0010" when "0101",
      "0000" when "0110",
      "0110" when "0111",
      "1010" when "1000",
      "0000" when "1001",
      "1000" when "1010",
      "0100" when "1011",
      "0001" when "1100",
      "0000" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0100" when "0000",
      "1000" when "0001",
      "0011" when "0010",
      "0010" when "0011",
      "0110" when "0100",
      "0101" when "0101",
      "0000" when "0110",
      "1001" when "0111",
      "0001" when "1000",
      "0000" when "1001",
      "1010" when "1010",
      "0111" when "1011",
      "1011" when "1100",
      "0000" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0101" when "0000",
      "0000" when "0001",
      "0001" when "0010",
      "0011" when "0011",
      "0000" when "0100",
      "0110" when "0101",
      "0100" when "0110",
      "0000" when "0111",
      "0000" when "1000",
      "0111" when "1001",
      "0000" when "1010",
      "1000" when "1011",
      "0000" when "1100",
      "0010" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0001" when "0000",
      "0000" when "0001",
      "0101" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0010" when "0101",
      "0111" when "0110",
      "0000" when "0111",
      "0100" when "1000",
      "0011" when "1001",
      "0000" when "1010",
      "1000" when "1011",
      "0000" when "1100",
      "0110" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "001" when "0000",
      "000" when "0001",
      "000" when "0010",
      "010" when "0011",
      "000" when "0100",
      "000" when "0101",
      "011" when "0110",
      "000" when "0111",
      "100" when "1000",
      "000" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "001" when "0000",
      "000" when "0001",
      "000" when "0010",
      "010" when "0011",
      "000" when "0100",
      "000" when "0101",
      "011" when "0110",
      "000" when "0111",
      "100" when "1000",
      "000" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "000" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "001" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "010" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 117 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      Y <= s116;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 137 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      Y <= s136;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 119 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      Y <= s118;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_120_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 120 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_120_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_120_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      Y <= s119;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_136_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 136 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_136_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_136_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      Y <= s135;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 124 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      Y <= s123;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_165_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 165 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_165_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_165_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
signal s160 : std_logic_vector(33 downto 0) := (others => '0');
signal s161 : std_logic_vector(33 downto 0) := (others => '0');
signal s162 : std_logic_vector(33 downto 0) := (others => '0');
signal s163 : std_logic_vector(33 downto 0) := (others => '0');
signal s164 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
      s160 <= "0000000000000000000000000000000000";
      s161 <= "0000000000000000000000000000000000";
      s162 <= "0000000000000000000000000000000000";
      s163 <= "0000000000000000000000000000000000";
      s164 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      s160 <= s159;
      s161 <= s160;
      s162 <= s161;
      s163 <= s162;
      s164 <= s163;
      Y <= s164;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_0 : in std_logic_vector(31 downto 0);
          R_U_0 : in std_logic_vector(31 downto 0);
          R_V_0 : in std_logic_vector(31 downto 0);
          R_W_0 : in std_logic_vector(31 downto 0);
          Inv_11_0 : out std_logic_vector(31 downto 0);
          Inv_12_0 : out std_logic_vector(31 downto 0);
          Inv_13_0 : out std_logic_vector(31 downto 0);
          Inv_21_0 : out std_logic_vector(31 downto 0);
          Inv_22_0 : out std_logic_vector(31 downto 0);
          Inv_23_0 : out std_logic_vector(31 downto 0);
          Inv_31_0 : out std_logic_vector(31 downto 0);
          Inv_32_0 : out std_logic_vector(31 downto 0);
          Inv_33_0 : out std_logic_vector(31 downto 0);
          Inv_41_0 : out std_logic_vector(31 downto 0);
          Inv_42_0 : out std_logic_vector(31 downto 0);
          Inv_43_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_14_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_14_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_7_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_12_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_9_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_133_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_120_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_136_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_165_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount141_out : std_logic_vector(3 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add31_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add31_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add31_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product431_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product431_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product481_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product491_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product491_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product611_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product611_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product811_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product811_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product811_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract1_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product45_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product45_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product45_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay145No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay154No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay154No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add31_4_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add31_4_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product811_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product811_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product45_4_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product45_4_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay154No8_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay154No7_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay151No4_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No4_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No1_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay156No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay145No3_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_12_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_13_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_21_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_22_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_23_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_31_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_32_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_33_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_41_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_42_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_43_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No5_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No120_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No121_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No7_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No9_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No4_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No124_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No122_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No8_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No123_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Add101_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Add101_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay116No4_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No39_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay42No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No6_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No11_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay41No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No4_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Add131_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Add131_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No9_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay118No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay130No5_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add31_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add31_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No83_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product112_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product112_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No82_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product431_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product431_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Product431_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Product431_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product491_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product491_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product512_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product512_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product512_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product512_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product512_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product512_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product512_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product512_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product611_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product611_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product611_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product611_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product811_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product811_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No12_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No24_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No13_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay72No3_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product45_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product45_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount141_instance: ModuloCounter_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount141_out);
Ldiff_UU_del_1_0_IEEE <= Ldiff_UU_del_1_0;
   Ldiff_UU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_0_out,
                 X => Ldiff_UU_del_1_0_IEEE);
Ldiff_UV_del_1_0_IEEE <= Ldiff_UV_del_1_0;
   Ldiff_UV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_0_out,
                 X => Ldiff_UV_del_1_0_IEEE);
Ldiff_UW_del_1_0_IEEE <= Ldiff_UW_del_1_0;
   Ldiff_UW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_0_out,
                 X => Ldiff_UW_del_1_0_IEEE);
Ldiff_VU_del_1_0_IEEE <= Ldiff_VU_del_1_0;
   Ldiff_VU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_0_out,
                 X => Ldiff_VU_del_1_0_IEEE);
Ldiff_VV_del_1_0_IEEE <= Ldiff_VV_del_1_0;
   Ldiff_VV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_0_out,
                 X => Ldiff_VV_del_1_0_IEEE);
Ldiff_VW_del_1_0_IEEE <= Ldiff_VW_del_1_0;
   Ldiff_VW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_0_out,
                 X => Ldiff_VW_del_1_0_IEEE);
Ldiff_WU_del_1_0_IEEE <= Ldiff_WU_del_1_0;
   Ldiff_WU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_0_out,
                 X => Ldiff_WU_del_1_0_IEEE);
Ldiff_WV_del_1_0_IEEE <= Ldiff_WV_del_1_0;
   Ldiff_WV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_0_out,
                 X => Ldiff_WV_del_1_0_IEEE);
Ldiff_WW_del_1_0_IEEE <= Ldiff_WW_del_1_0;
   Ldiff_WW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_0_out,
                 X => Ldiff_WW_del_1_0_IEEE);
R_U_0_IEEE <= R_U_0;
   R_U_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_0_out,
                 X => R_U_0_IEEE);
R_V_0_IEEE <= R_V_0;
   R_V_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_0_out,
                 X => R_V_0_IEEE);
R_W_0_IEEE <= R_W_0;
   R_W_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_0_out,
                 X => R_W_0_IEEE);

Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_0_impl_out,
                 X => Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast);

SharedReg554_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg161_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg161_out;
SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg255_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg255_out;
SharedReg134_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg134_out;
SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg41_out;
SharedReg162_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg162_out;
SharedReg75_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg75_out;
SharedReg553_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product108_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg162_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg75_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg161_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg255_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg134_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg274_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg274_out;
SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg21_out;
SharedReg570_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg35_out;
SharedReg352_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg352_out;
SharedReg353_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg353_out;
SharedReg278_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg278_out;
   MUX_Product108_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg274_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg35_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg278_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg21_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg34_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product108_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_1_impl_out,
                 X => Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast);

SharedReg50_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg50_out;
SharedReg80_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg80_out;
SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg168_out;
SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg47_out;
SharedReg115_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg115_out;
SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg168_out;
SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg47_out;
   MUX_Product108_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg50_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg80_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg115_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg47_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg554_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg168_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg373_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg395_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
SharedReg287_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg287_out;
SharedReg358_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg358_out;
SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg11_out;
SharedReg27_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg27_out;
SharedReg6_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg6_out;
   MUX_Product108_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg27_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg287_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg358_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product108_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_2_impl_out,
                 X => Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg142_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg142_out;
SharedReg415_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg57_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg57_out;
SharedReg59_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg59_out;
SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg54_out;
SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg118_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg118_out;
   MUX_Product108_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg142_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg54_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg118_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg415_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg57_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg59_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg6_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg319_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg380_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg325_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg325_out;
SharedReg397_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg397_out;
SharedReg20_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg16_out;
   MUX_Product108_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg6_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg325_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product108_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_3_impl_out,
                 X => Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg89_out;
SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg123_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg123_out;
SharedReg98_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg98_out;
SharedReg101_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg101_out;
SharedReg102_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg102_out;
SharedReg553_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg554_out;
SharedReg1_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product108_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg89_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg123_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg98_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg101_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg102_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_3_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_0_out,
                 Y => Delay1No6_out);

SharedReg560_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg6_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg327_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg387_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg332_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg332_out;
Delay154No8_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast <= Delay154No8_out;
SharedReg20_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product108_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg332_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay154No8_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_3_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product108_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_4_impl_out,
                 X => Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg427_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg427_out;
SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg128_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg128_out;
SharedReg67_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg184_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg184_out;
SharedReg104_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg104_out;
SharedReg428_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg428_out;
SharedReg131_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg131_out;
SharedReg553_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product108_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg554_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg427_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg128_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg184_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg104_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg428_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg131_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_4_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_0_out,
                 Y => Delay1No8_out);

SharedReg558_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg5_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg5_out;
SharedReg6_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg6_out;
SharedReg344_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg344_out;
SharedReg309_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg317_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg317_out;
SharedReg350_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg350_out;
SharedReg30_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product108_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg317_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg350_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg30_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg5_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg6_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg344_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product108_4_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product110_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_0_impl_out,
                 X => Delay1No10_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast);

SharedReg554_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg8_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg557_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg41_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg41_out;
SharedReg561_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg134_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg134_out;
SharedReg110_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg110_out;
SharedReg161_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg161_out;
SharedReg72_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg72_out;
SharedReg43_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg43_out;
SharedReg76_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg76_out;
SharedReg553_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product110_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg72_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg43_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg76_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg41_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg134_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg110_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg161_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_0_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_0_out,
                 Y => Delay1No10_out);

SharedReg371_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg371_out;
SharedReg13_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg27_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg6_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg406_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg365_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg365_out;
Delay151No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_14_cast <= Delay151No_out;
   MUX_Product110_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg371_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay151No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_0_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product110_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_1_impl_out,
                 X => Delay1No12_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg78_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg81_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
SharedReg553_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg8_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg557_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg47_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg47_out;
SharedReg561_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg137_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg137_out;
SharedReg77_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg77_out;
SharedReg195_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg195_out;
SharedReg114_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg114_out;
   MUX_Product110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg137_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg77_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg195_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg114_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg554_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg47_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_1_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_0_out,
                 Y => Delay1No12_out);

SharedReg29_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
SharedReg282_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg282_out;
Delay151No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast <= Delay151No1_out;
SharedReg288_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg288_out;
SharedReg13_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg5_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg5_out;
SharedReg372_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay151No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg288_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_1_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product110_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_2_impl_out,
                 X => Delay1No14_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg174_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg55_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg55_out;
SharedReg86_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg86_out;
SharedReg553_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg8_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg557_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg84_out;
SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg142_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg142_out;
   MUX_Product110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg142_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg84_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg55_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg86_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_2_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_0_out,
                 Y => Delay1No14_out);

SharedReg11_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg318_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg29_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg29_out;
SharedReg291_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg291_out;
Delay151No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast <= Delay151No2_out;
Delay154No7_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast <= Delay154No7_out;
SharedReg13_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
   MUX_Product110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg29_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay151No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay154No7_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_2_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product110_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_3_impl_out,
                 X => Delay1No16_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg123_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg89_out;
SharedReg148_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg148_out;
SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg61_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg61_out;
SharedReg65_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg65_out;
SharedReg553_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg554_out;
SharedReg8_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg557_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg123_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg148_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg61_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg65_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg554_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_3_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_0_out,
                 Y => Delay1No16_out);

SharedReg560_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg5_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg326_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg29_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg29_out;
SharedReg335_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg335_out;
Delay151No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast <= Delay151No3_out;
SharedReg316_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg316_out;
SharedReg13_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg21_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg29_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay151No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg316_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_3_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product110_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_4_impl_out,
                 X => Delay1No18_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg155_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg104_out;
SharedReg187_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg187_out;
SharedReg94_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg94_out;
SharedReg67_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg67_out;
SharedReg18_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg18_out;
SharedReg553_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product110_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg554_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg104_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg94_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg67_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg18_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_4_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_0_out,
                 Y => Delay1No18_out);

SharedReg558_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg26_out;
SharedReg22_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg571_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg343_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg29_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg402_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg402_out;
Delay151No4_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast <= Delay151No4_out;
SharedReg414_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg414_out;
SharedReg24_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg24_out;
SharedReg557_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product110_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay151No4_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg414_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg24_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg26_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product110_4_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product109_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_3_impl_out,
                 X => Delay1No20_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg422_out;
SharedReg61_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg61_out;
SharedReg89_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg89_out;
SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg422_out;
SharedReg149_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg149_out;
SharedReg40_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg40_out;
SharedReg31_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg554_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg554_out;
SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg422_out;
SharedReg557_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product109_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg61_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg89_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg422_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg149_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg40_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg554_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product109_3_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_0_out,
                 Y => Delay1No20_out);

SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg34_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg35_out;
SharedReg386_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg556_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg14_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg305_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg305_out;
SharedReg568_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg568_out;
SharedReg557_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product109_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg568_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg21_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg35_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg305_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product109_3_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product109_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_4_impl_out,
                 X => Delay1No22_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg128_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg561_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg94_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
SharedReg218_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg218_out;
SharedReg155_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg427_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg427_out;
SharedReg130_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg130_out;
SharedReg70_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg70_out;
SharedReg40_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg40_out;
SharedReg554_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg554_out;
SharedReg8_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg8_out;
SharedReg557_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product109_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg40_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg554_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg8_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg128_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg218_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg427_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg130_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg70_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product109_4_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_4_impl_0_out,
                 Y => Delay1No22_out);

SharedReg558_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg570_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg27_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg35_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg35_out;
SharedReg401_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg401_out;
SharedReg309_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg556_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg556_out;
SharedReg312_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg312_out;
SharedReg13_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product109_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg556_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg312_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg35_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg401_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product109_4_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_4_impl_1_out,
                 Y => Delay1No23_out);

Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast <= Delay1No24_out;
Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast <= Delay1No25_out;
   Product111_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_0_impl_out,
                 X => Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast);

SharedReg554_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg72_out;
SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg161_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg161_out;
SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg72_out;
SharedReg190_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg190_out;
SharedReg134_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg134_out;
SharedReg110_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg110_out;
SharedReg136_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg136_out;
SharedReg553_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product111_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg134_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg110_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg136_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg161_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg72_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg190_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_0_impl_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_0_out,
                 Y => Delay1No24_out);

SharedReg361_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg361_out;
SharedReg30_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg21_out;
SharedReg22_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg5_out;
SharedReg405_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg29_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg29_out;
SharedReg365_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg275_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg275_out;
   MUX_Product111_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg361_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg29_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg275_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg21_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg5_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_0_impl_1_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_1_out,
                 Y => Delay1No25_out);

Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No26_out;
Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No27_out;
   Product111_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_1_impl_out,
                 X => Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg261_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg138_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg138_out;
SharedReg553_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg77_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg77_out;
SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg168_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg168_out;
SharedReg114_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg114_out;
SharedReg231_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg231_out;
SharedReg372_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg138_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg168_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg114_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg231_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg554_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg77_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_1_impl_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_0_out,
                 Y => Delay1No26_out);

SharedReg394_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg359_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg359_out;
SharedReg297_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg297_out;
SharedReg30_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg11_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg11_out;
SharedReg571_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg571_out;
SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
   MUX_Product111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg571_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg359_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg297_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_1_impl_1_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_1_out,
                 Y => Delay1No27_out);

Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No28_out;
Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No29_out;
   Product111_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_2_impl_out,
                 X => Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg142_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg240_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg240_out;
SharedReg318_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg239_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg239_out;
SharedReg144_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg553_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg174_out;
SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg174_out;
   MUX_Product111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg240_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg174_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg239_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg144_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_2_impl_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_0_out,
                 Y => Delay1No28_out);

SharedReg33_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg571_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg571_out;
SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg379_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg291_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg398_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg398_out;
SharedReg340_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg340_out;
SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg15_out;
SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg26_out;
   MUX_Product111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg571_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg15_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg26_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg28_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg398_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg340_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_2_impl_1_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_1_out,
                 Y => Delay1No29_out);

Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast <= Delay1No30_out;
Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast <= Delay1No31_out;
   Product111_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_3_impl_out,
                 X => Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg148_out;
SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg123_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg123_out;
SharedReg246_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg246_out;
SharedReg326_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg210_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg210_out;
SharedReg125_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg125_out;
SharedReg553_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product111_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg148_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg123_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg246_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg210_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg125_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg554_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_3_impl_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_0_out,
                 Y => Delay1No30_out);

SharedReg560_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg33_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg33_out;
SharedReg571_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg571_out;
SharedReg28_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg386_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg335_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg306_out;
SharedReg342_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg342_out;
SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product111_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg33_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg571_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg342_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_3_impl_1_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_1_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Product111_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_4_impl_out,
                 X => Delay1No32_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg155_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg155_out;
SharedReg105_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg66_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg66_out;
SharedReg492_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg492_out;
SharedReg343_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg217_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg217_out;
SharedReg309_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg553_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg554_out;
SharedReg1_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product111_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg554_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg155_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg66_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg492_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg217_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_4_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_4_impl_0_out,
                 Y => Delay1No32_out);

SharedReg558_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg10_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg10_out;
SharedReg11_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg563_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg28_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg401_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg401_out;
SharedReg36_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg36_out;
SharedReg313_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg313_out;
Delay156No4_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast <= Delay156No4_out;
SharedReg13_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product111_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg313_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay156No4_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg15_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg10_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg563_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg401_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg36_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product111_4_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_4_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Product310_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_0_impl_out,
                 X => Delay1No34_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast);

SharedReg554_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg190_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg190_out;
SharedReg109_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg109_out;
SharedReg223_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg223_out;
SharedReg405_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg254_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg254_out;
SharedReg18_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg553_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product310_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg254_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg190_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg109_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg223_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_0_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_0_out,
                 Y => Delay1No34_out);

Delay156No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast <= Delay156No_out;
SharedReg24_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg557_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg26_out;
SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg28_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg352_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg352_out;
SharedReg353_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg353_out;
Delay156No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast <= Delay156No5_out;
   MUX_Product310_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay156No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay156No5_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg26_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_0_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Product310_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_1_impl_out,
                 X => Delay1No36_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast);

SharedReg230_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg18_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg553_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg168_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg168_out;
SharedReg195_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg195_out;
SharedReg137_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg461_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg461_out;
SharedReg12_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
   MUX_Product310_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg195_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg461_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg554_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg168_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_1_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_0_out,
                 Y => Delay1No36_out);

SharedReg281_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg281_out;
SharedReg395_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
Delay156No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast <= Delay156No6_out;
Delay156No1_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast <= Delay156No1_out;
SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg557_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg15_out;
SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg26_out;
SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg33_out;
SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
SharedReg372_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product310_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg281_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg26_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg33_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay156No6_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay156No1_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg15_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_1_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Product310_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_2_impl_out,
                 X => Delay1No38_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast);

SharedReg120_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg120_out;
SharedReg453_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg453_out;
SharedReg12_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg238_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg238_out;
SharedReg18_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg553_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg554_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg20_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg201_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg201_out;
SharedReg55_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg55_out;
   MUX_Product310_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg120_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg453_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg201_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg55_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg12_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg238_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_2_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_0_out,
                 Y => Delay1No38_out);

SharedReg22_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg318_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg290_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg290_out;
SharedReg380_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg299_out;
SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg299_out;
SharedReg24_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg557_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg10_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg10_out;
   MUX_Product310_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg10_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg290_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg299_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_2_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product310_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_3_impl_out,
                 X => Delay1No40_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg179_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg179_out;
SharedReg99_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg91_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg91_out;
SharedReg265_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg12_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg209_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg209_out;
SharedReg18_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg18_out;
SharedReg553_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg148_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg148_out;
SharedReg20_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product310_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg99_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg91_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg209_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg18_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg148_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_3_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_0_out,
                 Y => Delay1No40_out);

SharedReg560_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg10_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg326_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg334_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg334_out;
SharedReg387_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg342_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg342_out;
SharedReg567_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg24_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg557_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product310_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg10_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg334_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg342_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_3_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product310_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_4_impl_out,
                 X => Delay1No42_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg184_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg184_out;
SharedReg247_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg247_out;
SharedReg94_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg249_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg249_out;
SharedReg12_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg185_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg185_out;
SharedReg7_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg7_out;
SharedReg553_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg155_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg155_out;
SharedReg30_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg30_out;
SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product310_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg155_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg30_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg184_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg247_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg249_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg185_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg7_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_4_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_0_out,
                 Y => Delay1No42_out);

SharedReg558_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg33_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg33_out;
SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg343_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg308_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg402_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg402_out;
Delay156No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast <= Delay156No9_out;
SharedReg567_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg557_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product310_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay156No9_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg33_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product310_4_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Product610_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_0_impl_out,
                 X => Delay1No44_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast);

SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg161_out;
SharedReg42_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg42_out;
SharedReg134_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg134_out;
SharedReg458_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg458_out;
SharedReg12_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg222_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg222_out;
SharedReg365_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg553_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product610_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg222_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg161_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg42_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg134_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg458_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_0_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_0_out,
                 Y => Delay1No44_out);

SharedReg567_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg15_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg15_out;
SharedReg10_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg10_out;
SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg405_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg364_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg364_out;
SharedReg36_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg36_out;
SharedReg276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg276_out;
   MUX_Product610_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg364_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg36_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg557_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg15_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg10_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_0_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product610_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_1_impl_out,
                 X => Delay1No46_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast);

SharedReg197_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg197_out;
SharedReg282_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg553_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg137_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg137_out;
SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg195_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg195_out;
SharedReg48_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg116_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg116_out;
SharedReg451_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg451_out;
SharedReg280_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg280_out;
   MUX_Product610_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg197_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg116_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg451_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg280_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg195_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_1_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_0_out,
                 Y => Delay1No46_out);

SharedReg373_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg36_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg360_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg360_out;
SharedReg567_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg10_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg10_out;
SharedReg22_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg571_out;
SharedReg372_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product610_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg10_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg571_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg360_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_1_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product610_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_2_impl_out,
                 X => Delay1No48_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast);

SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg455_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg455_out;
SharedReg289_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg289_out;
SharedReg202_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg202_out;
SharedReg291_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg553_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg142_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg142_out;
SharedReg1_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg236_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg236_out;
SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg263_out;
   MUX_Product610_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg455_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg236_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg263_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg289_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg202_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg142_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_2_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_0_out,
                 Y => Delay1No48_out);

SharedReg11_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg571_out;
SharedReg318_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg319_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg36_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg399_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg399_out;
SharedReg567_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg557_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg558_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg16_out;
   MUX_Product610_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg571_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg16_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg399_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_2_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product610_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_3_impl_out,
                 X => Delay1No50_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast);

SharedReg123_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg208_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg243_out;
SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg489_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg489_out;
SharedReg333_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg333_out;
SharedReg181_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg181_out;
SharedReg335_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg553_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg179_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg179_out;
SharedReg1_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg14_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product610_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg489_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg333_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg181_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg179_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_3_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_0_out,
                 Y => Delay1No50_out);

SharedReg560_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg571_out;
SharedReg326_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg327_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg36_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg36_out;
Delay145No3_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast <= Delay145No3_out;
SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product610_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg571_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg36_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay145No3_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_3_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product610_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_4_impl_out,
                 X => Delay1No52_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg216_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg216_out;
SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg267_out;
SharedReg96_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg96_out;
SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg267_out;
SharedReg307_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg307_out;
SharedReg157_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg157_out;
SharedReg309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg553_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg184_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg184_out;
SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg14_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg14_out;
   MUX_Product610_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg184_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg14_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg216_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg96_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg267_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg307_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg157_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_4_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_0_out,
                 Y => Delay1No52_out);

SharedReg558_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg26_out;
SharedReg22_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg343_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg344_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg344_out;
SharedReg402_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg402_out;
SharedReg314_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg314_out;
SharedReg567_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg31_out;
   MUX_Product610_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg314_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg31_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg26_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg563_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg344_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product610_4_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product710_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_0_impl_out,
                 X => Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast);

SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg190_out;
SharedReg30_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg14_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg190_out;
SharedReg445_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg445_out;
SharedReg111_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg111_out;
SharedReg448_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg448_out;
SharedReg363_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg363_out;
SharedReg192_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg192_out;
SharedReg7_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg7_out;
SharedReg553_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product710_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg363_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg192_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg7_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg14_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg190_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg445_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg111_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg448_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_0_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_0_out,
                 Y => Delay1No54_out);

SharedReg567_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg571_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg405_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg406_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg353_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg353_out;
SharedReg279_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg279_out;
   MUX_Product710_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg279_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_0_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product710_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_1_impl_out,
                 X => Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast);

SharedReg450_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg450_out;
SharedReg7_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg553_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg168_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg168_out;
SharedReg30_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg229_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg229_out;
SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg449_out;
SharedReg258_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg258_out;
SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg449_out;
SharedReg12_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
   MUX_Product710_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg450_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg258_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg449_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg229_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_1_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_0_out,
                 Y => Delay1No56_out);

SharedReg373_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg395_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
SharedReg362_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg362_out;
SharedReg567_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg11_out;
SharedReg563_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
SharedReg372_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product710_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg362_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_1_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product710_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_2_impl_out,
                 X => Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast);

SharedReg144_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg144_out;
SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg263_out;
SharedReg12_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg454_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg454_out;
SharedReg7_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg553_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg174_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg174_out;
SharedReg30_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg14_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg118_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg118_out;
SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg263_out;
SharedReg453_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg453_out;
   MUX_Product710_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg144_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg263_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg453_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg12_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg454_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg174_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_2_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_0_out,
                 Y => Delay1No58_out);

SharedReg570_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg318_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg319_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg380_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg298_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg298_out;
SharedReg567_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg26_out;
   MUX_Product710_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg26_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg298_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_2_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product710_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_3_impl_out,
                 X => Delay1No60_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast);

SharedReg148_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg243_out;
SharedReg265_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg265_out;
SharedReg151_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg151_out;
SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg243_out;
SharedReg12_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg266_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg266_out;
SharedReg7_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg553_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg123_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg123_out;
SharedReg30_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg9_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product710_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg265_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg151_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg243_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg266_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg123_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_3_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_0_out,
                 Y => Delay1No60_out);

SharedReg560_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg570_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg326_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg327_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg387_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg341_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg341_out;
SharedReg567_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product710_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg26_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg341_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_3_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product710_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_4_impl_out,
                 X => Delay1No62_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg66_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg247_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg247_out;
SharedReg184_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg184_out;
SharedReg216_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg527_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg527_out;
SharedReg12_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg248_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg248_out;
SharedReg309_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg553_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg128_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg128_out;
SharedReg8_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg8_out;
SharedReg9_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg9_out;
   MUX_Product710_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg128_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg8_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg66_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg247_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg184_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg216_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg527_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg248_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_4_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_4_impl_0_out,
                 Y => Delay1No62_out);

SharedReg558_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg11_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg571_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg343_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg344_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg344_out;
SharedReg23_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg23_out;
SharedReg350_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg350_out;
SharedReg567_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Product710_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg350_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg344_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg23_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product710_4_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_4_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product810_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_0_impl_out,
                 X => Delay1No64_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg1_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg9_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg109_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg109_out;
SharedReg221_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg221_out;
SharedReg458_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg458_out;
SharedReg252_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg252_out;
SharedReg445_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg447_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg447_out;
SharedReg365_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg553_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product810_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg447_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg109_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg221_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg458_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg252_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_0_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_0_out,
                 Y => Delay1No64_out);

SharedReg567_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg26_out;
SharedReg11_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg405_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg406_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg353_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg353_out;
SharedReg277_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg277_out;
   MUX_Product810_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg277_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg26_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_0_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product810_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_1_impl_out,
                 X => Delay1No66_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast);

SharedReg441_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg441_out;
SharedReg282_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg553_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg1_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg9_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg114_out;
SharedReg258_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg258_out;
SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg461_out;
SharedReg138_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg138_out;
SharedReg463_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg463_out;
SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg461_out;
   MUX_Product810_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg441_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg138_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg463_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg461_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg114_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg258_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_1_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_0_out,
                 Y => Delay1No66_out);

SharedReg394_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg395_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
SharedReg286_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg26_out;
SharedReg570_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg571_out;
SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg564_out;
   MUX_Product810_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg26_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg571_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg564_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg286_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_1_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product810_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_2_impl_out,
                 X => Delay1No68_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast);

SharedReg482_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg482_out;
SharedReg485_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg485_out;
SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg453_out;
SharedReg509_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg509_out;
SharedReg291_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg553_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg118_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg118_out;
SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg9_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg142_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg142_out;
SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg453_out;
SharedReg201_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg201_out;
   MUX_Product810_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg482_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg485_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg142_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg201_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg453_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg509_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg118_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_2_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_0_out,
                 Y => Delay1No68_out);

SharedReg4_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg571_out;
SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg379_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg380_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg324_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg324_out;
SharedReg567_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg16_out;
   MUX_Product810_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg571_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg16_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg564_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg324_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_2_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product810_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_3_impl_out,
                 X => Delay1No70_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast);

SharedReg208_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg265_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg265_out;
SharedReg179_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg179_out;
SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg488_out;
SharedReg520_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg520_out;
SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg488_out;
SharedReg518_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg518_out;
SharedReg335_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg553_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg427_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg427_out;
SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product810_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg265_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg179_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg520_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg488_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg518_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg427_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_3_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_0_out,
                 Y => Delay1No70_out);

SharedReg560_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg4_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg571_out;
SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg564_out;
SharedReg386_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg387_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg339_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg339_out;
SharedReg567_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product810_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg571_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg564_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg339_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_3_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product810_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_4_impl_out,
                 X => Delay1No72_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg94_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg267_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg267_out;
SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg492_out;
SharedReg97_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg97_out;
SharedReg270_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg270_out;
SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg492_out;
SharedReg526_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg526_out;
SharedReg309_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg553_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg555_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg555_out;
SharedReg24_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg24_out;
SharedReg2_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
   MUX_Product810_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg555_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg24_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg94_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg267_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg97_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg270_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg492_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg526_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_4_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_0_out,
                 Y => Delay1No72_out);

SharedReg558_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg570_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg564_out;
SharedReg401_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg401_out;
SharedReg23_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg23_out;
SharedReg315_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg315_out;
SharedReg567_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Product810_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg315_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg564_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg401_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg23_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product810_4_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product910_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_0_impl_out,
                 X => Delay1No74_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast);

SharedReg433_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg433_out;
SharedReg8_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg2_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg134_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg134_out;
SharedReg252_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg252_out;
SharedReg221_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg221_out;
SharedReg136_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg136_out;
SharedReg467_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg467_out;
SharedReg466_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg466_out;
SharedReg500_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg500_out;
SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg553_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg553_out;
   MUX_Product910_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg433_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg466_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg500_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg134_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg252_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg221_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg136_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg467_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_0_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_0_out,
                 Y => Delay1No74_out);

SharedReg567_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg570_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg564_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg564_out;
SharedReg352_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg352_out;
SharedReg23_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg23_out;
SharedReg370_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg370_out;
   MUX_Product910_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg564_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg23_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg370_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_0_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product910_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_1_impl_out,
                 X => Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast);

SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg461_out;
SharedReg282_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg553_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg439_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg8_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg2_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg137_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg137_out;
SharedReg449_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg449_out;
SharedReg229_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg229_out;
SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg461_out;
SharedReg462_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg462_out;
SharedReg393_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg393_out;
   MUX_Product910_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg229_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg461_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg462_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg393_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg553_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg439_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg137_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg449_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_1_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_0_out,
                 Y => Delay1No76_out);

SharedReg281_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg281_out;
SharedReg23_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg285_out;
SharedReg567_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg16_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg4_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg571_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg571_out;
SharedReg17_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg17_out;
   MUX_Product910_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg281_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg571_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg17_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_1_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product910_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_2_impl_out,
                 X => Delay1No78_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast);

SharedReg455_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg455_out;
SharedReg484_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg484_out;
SharedReg378_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg378_out;
SharedReg453_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg453_out;
SharedReg291_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg553_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg422_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg422_out;
SharedReg8_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg2_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg201_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg201_out;
SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg482_out;
SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg482_out;
   MUX_Product910_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg455_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg484_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg201_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg482_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg378_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg453_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg422_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_2_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_0_out,
                 Y => Delay1No78_out);

SharedReg570_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg571_out;
SharedReg17_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
SharedReg290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg290_out;
SharedReg23_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg323_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg323_out;
SharedReg567_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg32_out;
   MUX_Product910_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg571_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg32_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg323_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_2_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product910_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_3_impl_out,
                 X => Delay1No80_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast);

SharedReg243_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg488_out;
SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg488_out;
SharedReg489_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg489_out;
SharedReg519_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg519_out;
SharedReg385_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg385_out;
SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg488_out;
SharedReg335_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg553_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg208_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg208_out;
SharedReg8_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg9_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product910_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg489_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg519_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg385_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg488_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg208_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_3_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_0_out,
                 Y => Delay1No80_out);

SharedReg560_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg570_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg571_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg571_out;
SharedReg17_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg334_out;
SharedReg23_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg331_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg331_out;
SharedReg567_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product910_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg571_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg17_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg331_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_3_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product910_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_4_impl_out,
                 X => Delay1No82_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg155_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg155_out;
SharedReg492_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg492_out;
SharedReg562_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg267_out;
SharedReg524_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg524_out;
SharedReg400_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg400_out;
SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg267_out;
SharedReg309_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg553_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg553_out;
SharedReg216_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg216_out;
SharedReg1_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg9_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg9_out;
   MUX_Product910_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg553_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg216_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg155_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg492_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg524_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg400_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg267_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_4_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_4_impl_0_out,
                 Y => Delay1No82_out);

SharedReg558_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg4_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg563_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg17_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg308_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg36_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg36_out;
SharedReg349_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg349_out;
SharedReg567_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg31_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg31_out;
   MUX_Product910_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg349_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg31_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg563_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg36_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product910_4_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_4_impl_1_out,
                 Y => Delay1No83_out);
   Inv_11_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_0_IEEE,
                 X => Delay1No84_out);
Inv_11_0 <= Inv_11_0_IEEE;

SharedReg41_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg47_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast <= SharedReg47_out;
SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg66_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast <= SharedReg66_out;
   MUX_Inv_11_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg66_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_11_0_0_LUT_out,
                 oMux => MUX_Inv_11_0_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_11_0_0_out,
                 Y => Delay1No84_out);
   Inv_12_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_0_IEEE,
                 X => Delay1No85_out);
Inv_12_0 <= Inv_12_0_IEEE;

SharedReg72_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg77_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg84_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg89_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast <= SharedReg89_out;
SharedReg94_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
   MUX_Inv_12_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg84_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg89_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_12_0_0_LUT_out,
                 oMux => MUX_Inv_12_0_0_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_12_0_0_out,
                 Y => Delay1No85_out);
   Inv_13_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_0_IEEE,
                 X => Delay1No86_out);
Inv_13_0 <= Inv_13_0_IEEE;

SharedReg72_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg77_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg84_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg60_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg66_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast <= SharedReg66_out;
   MUX_Inv_13_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg84_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg66_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_13_0_0_LUT_out,
                 oMux => MUX_Inv_13_0_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_13_0_0_out,
                 Y => Delay1No86_out);
   Inv_21_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_0_IEEE,
                 X => Delay1No87_out);
Inv_21_0 <= Inv_21_0_IEEE;

SharedReg134_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg137_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast <= SharedReg148_out;
SharedReg155_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
   MUX_Inv_21_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_21_0_0_LUT_out,
                 oMux => MUX_Inv_21_0_0_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_21_0_0_out,
                 Y => Delay1No87_out);
   Inv_22_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_0_IEEE,
                 X => Delay1No88_out);
Inv_22_0 <= Inv_22_0_IEEE;

SharedReg109_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast <= SharedReg109_out;
SharedReg114_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast <= SharedReg114_out;
SharedReg118_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast <= SharedReg89_out;
SharedReg94_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
   MUX_Inv_22_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg109_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg118_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg89_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_22_0_0_LUT_out,
                 oMux => MUX_Inv_22_0_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_22_0_0_out,
                 Y => Delay1No88_out);
   Inv_23_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_0_IEEE,
                 X => Delay1No89_out);
Inv_23_0 <= Inv_23_0_IEEE;

SharedReg134_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg123_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast <= SharedReg123_out;
SharedReg128_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast <= SharedReg128_out;
   MUX_Inv_23_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg123_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg128_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_23_0_0_LUT_out,
                 oMux => MUX_Inv_23_0_0_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_23_0_0_out,
                 Y => Delay1No89_out);
   Inv_31_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_0_IEEE,
                 X => Delay1No90_out);
Inv_31_0 <= Inv_31_0_IEEE;

SharedReg161_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg168_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast <= SharedReg168_out;
SharedReg174_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg179_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast <= SharedReg179_out;
SharedReg184_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast <= SharedReg184_out;
   MUX_Inv_31_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg168_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg179_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg184_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_31_0_0_LUT_out,
                 oMux => MUX_Inv_31_0_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_31_0_0_out,
                 Y => Delay1No90_out);
   Inv_32_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_0_IEEE,
                 X => Delay1No91_out);
Inv_32_0 <= Inv_32_0_IEEE;

SharedReg190_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast <= SharedReg190_out;
SharedReg195_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast <= SharedReg195_out;
SharedReg201_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast <= SharedReg201_out;
SharedReg208_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast <= SharedReg208_out;
SharedReg216_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast <= SharedReg216_out;
   MUX_Inv_32_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg190_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg201_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg208_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg216_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_32_0_0_LUT_out,
                 oMux => MUX_Inv_32_0_0_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_32_0_0_out,
                 Y => Delay1No91_out);
   Inv_33_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_0_IEEE,
                 X => Delay1No92_out);
Inv_33_0 <= Inv_33_0_IEEE;

SharedReg221_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg229_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast <= SharedReg229_out;
SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg247_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast <= SharedReg247_out;
   MUX_Inv_33_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg236_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg247_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_33_0_0_LUT_out,
                 oMux => MUX_Inv_33_0_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_33_0_0_out,
                 Y => Delay1No92_out);
   Inv_41_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_0_IEEE,
                 X => Delay1No93_out);
Inv_41_0 <= Inv_41_0_IEEE;

SharedReg252_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg258_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast <= SharedReg258_out;
SharedReg263_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg265_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg267_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast <= SharedReg267_out;
   MUX_Inv_41_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg258_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg263_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_41_0_0_LUT_out,
                 oMux => MUX_Inv_41_0_0_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_41_0_0_out,
                 Y => Delay1No93_out);
   Inv_42_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_0_IEEE,
                 X => Delay1No94_out);
Inv_42_0 <= Inv_42_0_IEEE;

SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg47_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast <= SharedReg47_out;
SharedReg54_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg98_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg104_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
   MUX_Inv_42_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_42_0_0_LUT_out,
                 oMux => MUX_Inv_42_0_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_42_0_0_out,
                 Y => Delay1No94_out);
   Inv_43_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_0_IEEE,
                 X => Delay1No95_out);
Inv_43_0 <= Inv_43_0_IEEE;

SharedReg109_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast <= SharedReg109_out;
SharedReg114_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast <= SharedReg114_out;
SharedReg118_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg123_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast <= SharedReg123_out;
SharedReg128_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast <= SharedReg128_out;
   MUX_Inv_43_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg109_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg118_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg123_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg128_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Inv_43_0_0_LUT_out,
                 oMux => MUX_Inv_43_0_0_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_43_0_0_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_0_impl_out,
                 X => Delay1No96_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast);

Delay16No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast <= Delay16No_out;
SharedReg190_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg190_out;
Delay22No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast <= Delay22No_out;
Delay22No5_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast <= Delay22No5_out;
SharedReg225_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg225_out;
SharedReg504_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg504_out;
SharedReg471_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg471_out;
SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg45_out;
SharedReg164_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg164_out;
SharedReg112_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg112_out;
SharedReg252_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg252_out;
SharedReg46_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg221_out;
SharedReg446_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg446_out;
   MUX_Add30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay16No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg190_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg252_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg446_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay22No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay22No5_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg225_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg504_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg471_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg45_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg164_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg112_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_0_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_0_out,
                 Y => Delay1No96_out);

Delay2No120_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast <= Delay2No120_out;
SharedReg252_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg363_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg363_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg547_out;
SharedReg405_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
SharedReg271_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg271_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg547_out;
SharedReg445_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg445_out;
SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg547_out;
SharedReg191_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg191_out;
SharedReg72_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg72_out;
   MUX_Add30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No120_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg445_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg191_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg72_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg363_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg271_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg547_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_0_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_1_impl_out,
                 X => Delay1No98_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg53_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg195_out;
SharedReg259_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg259_out;
Delay16No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast <= Delay16No1_out;
SharedReg168_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg168_out;
Delay22No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast <= Delay22No1_out;
Delay22No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast <= Delay22No6_out;
SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg195_out;
SharedReg_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
Delay116No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast <= Delay116No1_out;
SharedReg83_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg83_out;
SharedReg233_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg233_out;
SharedReg77_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg77_out;
Delay13No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast <= Delay13No6_out;
   MUX_Add30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg83_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg233_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg77_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay13No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg259_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay16No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg168_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay22No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay22No6_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg195_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay116No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_1_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_0_out,
                 Y => Delay1No98_out);

SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg548_out;
SharedReg196_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg196_out;
SharedReg47_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg47_out;
Delay2No121_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast <= Delay2No121_out;
SharedReg229_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg229_out;
SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg548_out;
SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg372_out;
SharedReg283_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg283_out;
SharedReg473_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg473_out;
SharedReg377_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg377_out;
SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg548_out;
SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg372_out;
SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg114_out;
SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg548_out;
   MUX_Add30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg196_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg114_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg47_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No121_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg229_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg548_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg372_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg283_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg473_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg377_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_1_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_2_impl_out,
                 X => Delay1No100_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast);

SharedReg145_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg121_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg201_out;
SharedReg173_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg173_out;
Delay45No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast <= Delay45No1_out;
Delay42No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast <= Delay42No1_out;
SharedReg444_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg444_out;
SharedReg174_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg174_out;
SharedReg420_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg420_out;
SharedReg147_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg147_out;
SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg201_out;
SharedReg_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg_out;
Delay116No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast <= Delay116No2_out;
Delay11No7_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast <= Delay11No7_out;
   MUX_Add30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay116No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay11No7_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg201_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg173_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay45No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay42No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg444_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg174_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg420_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg147_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_2_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_0_out,
                 Y => Delay1No100_out);

SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg549_out;
SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg549_out;
SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg548_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg548_out;
SharedReg373_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg373_out;
SharedReg396_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg396_out;
SharedReg375_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg375_out;
SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg549_out;
SharedReg378_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg378_out;
SharedReg321_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg321_out;
SharedReg507_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg507_out;
SharedReg322_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg322_out;
SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg549_out;
   MUX_Add30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg321_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg507_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg322_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg548_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg373_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg375_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg236_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg549_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg378_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_2_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add30_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_3_impl_out,
                 X => Delay1No102_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast);

SharedReg538_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg538_out;
SharedReg490_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg490_out;
SharedReg423_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg423_out;
SharedReg84_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg84_out;
SharedReg486_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg486_out;
SharedReg512_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg512_out;
SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg54_out;
Delay45No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast <= Delay45No2_out;
Delay42No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast <= Delay42No2_out;
SharedReg515_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg515_out;
SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg179_out;
SharedReg424_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg424_out;
SharedReg154_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg154_out;
SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg179_out;
   MUX_Add30_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg538_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg490_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg424_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg154_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg179_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg423_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg84_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg486_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg512_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg54_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay45No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay42No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg515_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_3_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_0_out,
                 Y => Delay1No102_out);

SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg551_out;
SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg326_out;
SharedReg300_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg300_out;
SharedReg118_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg118_out;
SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg549_out;
SharedReg319_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg319_out;
SharedReg56_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg56_out;
SharedReg379_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg379_out;
SharedReg382_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg382_out;
SharedReg381_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg381_out;
SharedReg243_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg243_out;
SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg326_out;
SharedReg329_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg329_out;
   MUX_Add30_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg243_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg326_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg329_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg300_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg118_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg549_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg319_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg56_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg379_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg382_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg381_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_3_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add30_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_4_impl_out,
                 X => Delay1No104_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast);

Delay22No9_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast <= Delay22No9_out;
SharedReg219_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg219_out;
SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg_out;
SharedReg528_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg528_out;
SharedReg107_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg107_out;
SharedReg159_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg159_out;
SharedReg89_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg89_out;
SharedReg216_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg216_out;
SharedReg430_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg430_out;
SharedReg153_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg153_out;
SharedReg268_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg268_out;
Delay16No4_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast <= Delay16No4_out;
SharedReg184_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg184_out;
SharedReg104_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg104_out;
   MUX_Add30_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay22No9_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg219_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg268_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay16No4_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg184_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg104_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg528_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg107_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg159_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg89_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg216_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg430_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg153_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_4_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_0_out,
                 Y => Delay1No104_out);

SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg551_out;
SharedReg492_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg492_out;
SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
SharedReg385_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg385_out;
SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg550_out;
SharedReg123_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg247_out;
SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg550_out;
SharedReg549_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg549_out;
SharedReg104_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg104_out;
Delay2No124_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast <= Delay2No124_out;
SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg247_out;
SharedReg129_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg129_out;
   MUX_Add30_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg551_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg104_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay2No124_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg129_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg492_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg385_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg247_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg550_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg549_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add30_4_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add110_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_2_impl_out,
                 X => Delay1No106_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg206_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg54_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg54_out;
SharedReg88_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg419_out;
SharedReg174_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg174_out;
SharedReg237_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg237_out;
Delay16No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast <= Delay16No2_out;
SharedReg263_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg263_out;
SharedReg84_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg84_out;
SharedReg242_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg242_out;
Delay118No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast <= Delay118No2_out;
SharedReg19_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg19_out;
Delay130No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast <= Delay130No7_out;
SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg511_out;
   MUX_Add110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay118No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg19_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay130No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg88_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg174_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg237_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay16No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg263_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg84_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg242_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add110_2_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_0_out,
                 Y => Delay1No106_out);

SharedReg318_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg318_out;
SharedReg84_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg84_out;
SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg549_out;
SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg549_out;
SharedReg175_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
Delay2No122_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast <= Delay2No122_out;
SharedReg85_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg85_out;
SharedReg119_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg119_out;
SharedReg548_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg548_out;
SharedReg304_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg304_out;
SharedReg422_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg422_out;
SharedReg294_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg294_out;
SharedReg378_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg378_out;
   MUX_Add110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg318_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg304_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg422_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg294_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg378_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg549_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay2No122_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg85_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg119_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg548_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add110_2_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Add110_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_3_impl_out,
                 X => Delay1No108_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg19_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg19_out;
Delay130No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast <= Delay130No8_out;
SharedReg535_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg535_out;
SharedReg214_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg214_out;
SharedReg98_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg98_out;
SharedReg93_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg93_out;
SharedReg103_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg103_out;
SharedReg265_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg265_out;
SharedReg123_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg123_out;
SharedReg100_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg100_out;
SharedReg522_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg522_out;
SharedReg427_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg427_out;
Delay88No3_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast <= Delay88No3_out;
SharedReg491_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg491_out;
   MUX_Add110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay130No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg522_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg427_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay88No3_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg491_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg535_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg214_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg98_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg93_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg103_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg265_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg123_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg100_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add110_3_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_0_out,
                 Y => Delay1No108_out);

SharedReg427_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg336_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg336_out;
SharedReg326_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg326_out;
SharedReg333_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg333_out;
SharedReg60_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg551_out;
SharedReg549_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg549_out;
SharedReg213_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg213_out;
SharedReg338_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg338_out;
SharedReg98_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg98_out;
SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg551_out;
SharedReg522_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg522_out;
SharedReg387_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg387_out;
SharedReg385_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg385_out;
   MUX_Add110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg522_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg387_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg385_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg326_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg551_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg549_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg213_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg338_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg98_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add110_3_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Add101_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_3_impl_out,
                 X => Delay1No110_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
Delay116No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast <= Delay116No3_out;
Delay11No8_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast <= Delay11No8_out;
SharedReg152_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg126_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg126_out;
SharedReg208_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg208_out;
SharedReg146_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg146_out;
SharedReg179_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg179_out;
SharedReg244_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg244_out;
Delay16No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast <= Delay16No3_out;
SharedReg265_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg265_out;
SharedReg89_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg215_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg215_out;
Delay118No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_14_cast <= Delay118No3_out;
   MUX_Add101_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay116No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg265_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg215_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay118No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay11No8_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg152_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg208_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg146_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg179_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg244_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay16No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add101_3_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_3_impl_0_out,
                 Y => Delay1No110_out);

SharedReg532_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg532_out;
SharedReg337_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg337_out;
SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg551_out;
SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg551_out;
SharedReg243_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg243_out;
SharedReg548_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg548_out;
SharedReg180_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg180_out;
SharedReg60_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
Delay2No123_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast <= Delay2No123_out;
SharedReg90_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg90_out;
SharedReg124_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg124_out;
SharedReg549_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg549_out;
SharedReg391_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg391_out;
   MUX_Add101_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg532_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg90_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg124_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg549_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg391_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg551_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg243_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg548_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg180_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay2No123_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add101_3_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_3_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Add101_4_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Add101_4_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Add101_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_4_impl_out,
                 X => Delay1No112_out_to_Add101_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Add101_4_impl_parent_implementedSystem_port_1_cast);

SharedReg220_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg184_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg184_out;
SharedReg19_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg19_out;
Delay116No4_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_4_cast <= Delay116No4_out;
SharedReg108_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg108_out;
SharedReg251_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg251_out;
SharedReg71_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg71_out;
SharedReg132_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg132_out;
SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg216_out;
SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg216_out;
SharedReg94_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg94_out;
SharedReg68_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg68_out;
SharedReg267_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg267_out;
SharedReg524_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg524_out;
   MUX_Add101_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg94_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg68_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg267_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg524_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg19_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay116No4_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg108_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg251_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg71_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg132_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg216_out_to_MUX_Add101_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add101_4_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_4_impl_0_out,
                 Y => Delay1No112_out);

SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg550_out;
SharedReg403_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg524_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg524_out;
Delay12No39_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_4_cast <= Delay12No39_out;
SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg550_out;
SharedReg343_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg343_out;
SharedReg551_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg551_out;
SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg247_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg247_out;
SharedReg156_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg156_out;
SharedReg311_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg311_out;
SharedReg104_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg104_out;
SharedReg95_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg95_out;
SharedReg495_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg495_out;
   MUX_Add101_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg311_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg104_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg95_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg495_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg524_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay12No39_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg343_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg551_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg247_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg156_out_to_MUX_Add101_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add101_4_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_4_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Add111_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_1_impl_out,
                 X => Delay1No114_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg167_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg167_out;
Delay45No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast <= Delay45No_out;
Delay42No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast <= Delay42No_out;
SharedReg505_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg505_out;
SharedReg460_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg460_out;
SharedReg37_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg37_out;
SharedReg438_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg438_out;
SharedReg199_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg199_out;
SharedReg443_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg443_out;
SharedReg465_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg465_out;
SharedReg437_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg437_out;
SharedReg139_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg139_out;
SharedReg117_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg117_out;
SharedReg229_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg229_out;
   MUX_Add111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay45No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg437_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg139_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg117_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg229_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay42No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg505_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg460_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg37_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg438_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg199_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg443_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg465_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add111_1_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_0_out,
                 Y => Delay1No114_out);

SharedReg547_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg547_out;
SharedReg406_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg406_out;
SharedReg354_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg354_out;
SharedReg408_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg408_out;
SharedReg405_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg405_out;
SharedReg433_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg433_out;
SharedReg351_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg351_out;
SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg548_out;
SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg548_out;
SharedReg393_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg393_out;
SharedReg280_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg280_out;
SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg548_out;
SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg548_out;
SharedReg258_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg258_out;
   MUX_Add111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg547_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg406_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg280_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg258_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg354_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg408_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg405_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg433_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg351_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg548_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg393_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add111_1_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Add121_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_0_impl_out,
                 X => Delay1No116_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg445_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg72_out;
SharedReg226_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg226_out;
SharedReg190_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg190_out;
SharedReg_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
SharedReg506_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg506_out;
Delay11No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast <= Delay11No5_out;
SharedReg257_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg257_out;
SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg72_out;
Delay13No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast <= Delay13No5_out;
SharedReg252_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg252_out;
SharedReg458_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg458_out;
SharedReg134_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg134_out;
   MUX_Add121_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay13No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg252_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg458_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg134_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg226_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg190_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg506_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay11No5_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg257_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg72_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_0_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_0_out,
                 Y => Delay1No116_out);

SharedReg41_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg110_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg135_out;
SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg547_out;
SharedReg366_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg366_out;
SharedReg466_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg466_out;
SharedReg409_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg409_out;
SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg547_out;
SharedReg363_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg363_out;
SharedReg109_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg109_out;
SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg547_out;
SharedReg445_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg445_out;
SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg256_out;
SharedReg273_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg273_out;
   MUX_Add121_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg445_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg273_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg135_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg366_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg466_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg409_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg547_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg363_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg109_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_0_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Add121_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_1_impl_out,
                 X => Delay1No118_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast);

SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg449_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg449_out;
SharedReg114_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg49_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg49_out;
SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg258_out;
SharedReg77_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg77_out;
SharedReg234_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg234_out;
Delay118No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast <= Delay118No1_out;
SharedReg19_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg19_out;
Delay130No6_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast <= Delay130No6_out;
SharedReg478_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg478_out;
Delay82No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast <= Delay82No1_out;
SharedReg480_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg480_out;
SharedReg481_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg481_out;
   MUX_Add121_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg449_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg478_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay82No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg480_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg481_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg114_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg49_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg258_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg77_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg234_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay118No1_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg19_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay130No6_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_1_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_0_out,
                 Y => Delay1No118_out);

SharedReg449_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg449_out;
Delay18No11_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast <= Delay18No11_out;
SharedReg357_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg357_out;
SharedReg433_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg433_out;
SharedReg78_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg78_out;
SharedReg115_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg115_out;
SharedReg547_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg547_out;
SharedReg295_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg295_out;
SharedReg439_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg439_out;
SharedReg284_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg284_out;
SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg393_out;
SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg393_out;
SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg393_out;
SharedReg351_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg351_out;
   MUX_Add121_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg449_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay18No11_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg393_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg351_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg357_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg433_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg78_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg115_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg547_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg295_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg439_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg284_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_1_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Add121_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_2_impl_out,
                 X => Delay1No120_out_to_Add121_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Add121_2_impl_parent_implementedSystem_port_1_cast);

SharedReg426_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg426_out;
SharedReg513_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg513_out;
SharedReg514_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg514_out;
SharedReg236_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg263_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg263_out;
SharedReg118_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg417_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg417_out;
SharedReg487_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg487_out;
SharedReg422_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg422_out;
Delay88No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast <= Delay88No2_out;
SharedReg457_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg457_out;
SharedReg37_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg37_out;
Delay41No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast <= Delay41No2_out;
SharedReg213_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg213_out;
   MUX_Add121_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg426_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg513_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg457_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg37_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay41No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg213_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg514_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg263_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg118_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg417_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg487_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg422_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay88No2_out_to_MUX_Add121_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_2_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_2_impl_0_out,
                 Y => Delay1No120_out);

SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg378_out;
SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg378_out;
SharedReg393_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg393_out;
SharedReg263_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg263_out;
SharedReg241_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg241_out;
SharedReg296_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg296_out;
SharedReg415_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg415_out;
SharedReg549_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg549_out;
SharedReg487_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg487_out;
SharedReg380_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg380_out;
SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg300_out;
SharedReg98_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg98_out;
SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg300_out;
SharedReg551_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg551_out;
   MUX_Add121_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg378_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg300_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg551_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg393_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg263_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg241_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg296_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg415_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg549_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg487_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg380_out_to_MUX_Add121_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_2_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_2_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Add121_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_3_impl_out,
                 X => Delay1No122_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast);

SharedReg37_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg431_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg431_out;
SharedReg530_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg530_out;
SharedReg432_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg432_out;
SharedReg537_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg537_out;
Delay73No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast <= Delay73No3_out;
SharedReg243_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg243_out;
SharedReg521_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg521_out;
SharedReg536_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg536_out;
SharedReg60_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg60_out;
Delay45No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast <= Delay45No3_out;
SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg523_out;
SharedReg539_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg539_out;
Delay22No4_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast <= Delay22No4_out;
   MUX_Add121_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg431_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay45No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg523_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg539_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay22No4_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg530_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg432_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg537_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay73No3_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg243_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg521_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg536_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg60_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_3_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_0_out,
                 Y => Delay1No122_out);

SharedReg104_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg385_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg385_out;
SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg550_out;
SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg300_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
SharedReg265_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg265_out;
SharedReg551_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg327_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg327_out;
SharedReg62_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg386_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg386_out;
SharedReg389_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg389_out;
SharedReg388_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg388_out;
SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg550_out;
   MUX_Add121_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg385_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg386_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg389_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg388_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg550_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg265_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg327_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add121_3_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Add131_2_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Add131_2_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Add131_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_2_impl_out,
                 X => Delay1No124_out_to_Add131_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Add131_2_impl_parent_implementedSystem_port_1_cast);

SharedReg114_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg476_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg476_out;
SharedReg479_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg479_out;
SharedReg47_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg47_out;
SharedReg477_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg477_out;
SharedReg439_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg439_out;
Delay88No1_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_7_cast <= Delay88No1_out;
SharedReg452_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg452_out;
SharedReg37_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg37_out;
SharedReg421_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg421_out;
SharedReg205_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg205_out;
SharedReg425_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg425_out;
SharedReg456_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg456_out;
SharedReg442_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg442_out;
   MUX_Add131_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg476_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg205_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg425_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg456_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg442_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg479_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg47_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg477_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg439_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay88No1_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg452_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg37_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg421_out_to_MUX_Add131_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add131_2_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_2_impl_0_out,
                 Y => Delay1No124_out);

SharedReg137_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg548_out;
SharedReg373_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg373_out;
SharedReg79_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg79_out;
SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg464_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg464_out;
SharedReg374_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg374_out;
SharedReg393_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg393_out;
SharedReg415_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg415_out;
SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg289_out;
SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg549_out;
SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg549_out;
SharedReg378_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg378_out;
SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg289_out;
   MUX_Add131_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg549_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg378_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg373_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg79_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg464_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg374_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg393_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg415_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg289_out_to_MUX_Add131_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add131_2_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_2_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Add18_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_4_impl_out,
                 X => Delay1No126_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast);

Delay88No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast <= Delay88No4_out;
Delay118No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast <= Delay118No4_out;
SharedReg37_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg37_out;
Delay130No9_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast <= Delay130No9_out;
SharedReg544_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg544_out;
Delay82No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast <= Delay82No4_out;
SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg66_out;
SharedReg497_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg497_out;
SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg66_out;
SharedReg492_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg492_out;
SharedReg496_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg496_out;
SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg66_out;
SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg543_out;
SharedReg529_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg529_out;
   MUX_Add18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay88No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay118No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg496_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg529_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg37_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay130No9_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg544_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay82No4_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg497_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg66_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg492_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_4_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_0_out,
                 Y => Delay1No126_out);

SharedReg402_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg402_out;
SharedReg413_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg413_out;
SharedReg540_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg540_out;
SharedReg347_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg343_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg343_out;
SharedReg400_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg94_out;
SharedReg385_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg385_out;
SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg94_out;
SharedReg250_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg250_out;
SharedReg401_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg401_out;
SharedReg96_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg96_out;
SharedReg551_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg551_out;
SharedReg412_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg412_out;
   MUX_Add18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg402_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg413_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg401_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg96_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg551_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg412_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg540_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg385_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg94_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg250_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_4_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Add24_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_0_impl_out,
                 X => Delay1No128_out_to_Add24_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Add24_0_impl_parent_implementedSystem_port_1_cast);

SharedReg72_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg502_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg502_out;
SharedReg498_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg498_out;
Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast <= Delay88No_out;
Delay118No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast <= Delay118No_out;
SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg19_out;
Delay130No5_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast <= Delay130No5_out;
SharedReg470_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg470_out;
Delay82No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast <= Delay82No_out;
SharedReg503_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg503_out;
Delay73No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast <= Delay73No_out;
SharedReg109_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg109_out;
SharedReg468_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg468_out;
SharedReg472_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg472_out;
   MUX_Add24_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg502_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay73No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg109_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg468_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg472_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg498_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay88No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay118No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg19_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay130No5_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg470_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay82No_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg503_out_to_MUX_Add24_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add24_0_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_0_impl_0_out,
                 Y => Delay1No128_out);

SharedReg111_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg547_out;
SharedReg469_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg407_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg356_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg356_out;
SharedReg498_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg498_out;
SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg368_out;
SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg405_out;
SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg405_out;
SharedReg351_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg351_out;
SharedReg271_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg271_out;
SharedReg134_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg134_out;
SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg547_out;
SharedReg406_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg406_out;
   MUX_Add24_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg271_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg134_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg547_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg406_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg469_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg356_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg498_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg368_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg405_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg351_out_to_MUX_Add24_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add24_0_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_0_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add31_4_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add31_4_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add31_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add31_4_impl_out,
                 X => Delay1No130_out_to_Add31_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add31_4_impl_parent_implementedSystem_port_1_cast);

SharedReg133_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg494_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg494_out;
SharedReg531_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg531_out;
SharedReg546_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg546_out;
Delay45No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_5_cast <= Delay45No4_out;
SharedReg545_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg545_out;
Delay34No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_7_cast <= Delay34No4_out;
   MUX_Add31_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg494_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg531_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg546_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay45No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg545_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay34No4_out_to_MUX_Add31_4_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_Add31_4_impl_0_LUT_out,
                 oMux => MUX_Add31_4_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add31_4_impl_0_out,
                 Y => Delay1No130_out);

SharedReg551_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg551_out;
SharedReg550_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg550_out;
SharedReg403_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg403_out;
SharedReg400_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg410_out;
SharedReg411_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg411_out;
SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
   MUX_Add31_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg551_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg550_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg403_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg411_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Add31_4_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => MUX_Add31_4_impl_1_LUT_out,
                 oMux => MUX_Add31_4_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add31_4_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product112_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_2_impl_out,
                 X => Delay1No132_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast);

SharedReg85_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg118_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg439_out;
SharedReg176_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg176_out;
SharedReg40_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg439_out;
SharedReg461_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg461_out;
SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg450_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg450_out;
SharedReg174_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg174_out;
SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg415_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg415_out;
   MUX_Product112_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg450_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg174_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg415_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg176_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg439_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg461_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_2_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_0_out,
                 Y => Delay1No132_out);

SharedReg11_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg34_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg35_out;
SharedReg379_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg556_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg569_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg569_out;
SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
   MUX_Product112_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg569_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg35_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg568_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_2_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product112_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_3_impl_out,
                 X => Delay1No134_out_to_Product112_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product112_3_impl_parent_implementedSystem_port_1_cast);

SharedReg179_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg6_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
Delay7No83_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast <= Delay7No83_out;
SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg507_out;
SharedReg263_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg263_out;
SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg482_out;
SharedReg39_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg39_out;
SharedReg9_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg507_out;
SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg482_out;
SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg454_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg454_out;
   MUX_Product112_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg454_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg6_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No83_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg507_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg263_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg482_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg39_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product112_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_3_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_3_impl_0_out,
                 Y => Delay1No134_out);

SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg378_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg378_out;
SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg572_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg31_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg569_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg569_out;
   MUX_Product112_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg568_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg569_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg378_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg572_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg573_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product112_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_3_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_3_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product112_4_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product112_4_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product112_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_4_impl_out,
                 X => Delay1No136_out_to_Product112_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product112_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg266_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg561_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg427_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg427_out;
SharedReg6_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg128_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg128_out;
SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg532_out;
SharedReg265_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg265_out;
SharedReg106_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg106_out;
SharedReg39_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg39_out;
SharedReg31_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg1_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg532_out;
   MUX_Product112_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg39_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg266_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg427_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg128_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg532_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg265_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg106_out_to_MUX_Product112_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_4_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_4_impl_0_out,
                 Y => Delay1No136_out);

SharedReg558_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg569_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg561_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg21_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg385_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg385_out;
SharedReg34_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg34_out;
SharedReg572_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg573_out;
SharedReg402_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg402_out;
SharedReg556_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg556_out;
SharedReg14_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg20_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg568_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
   MUX_Product112_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg556_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg385_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg34_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg572_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg573_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Product112_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product112_4_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_4_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product102_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_1_impl_out,
                 X => Delay1No138_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast);

SharedReg169_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg40_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg31_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg498_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg498_out;
SharedReg458_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg458_out;
SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg433_out;
SharedReg447_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg447_out;
SharedReg501_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg6_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg262_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg262_out;
SharedReg137_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg137_out;
SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg433_out;
   MUX_Product102_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg262_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg137_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg498_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg458_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg433_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg447_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product102_1_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_0_out,
                 Y => Delay1No138_out);

SharedReg394_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg556_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg14_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg558_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg351_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg351_out;
SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg34_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg34_out;
SharedReg35_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg35_out;
   MUX_Product102_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg351_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg34_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg35_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg14_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg568_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg569_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product102_1_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product102_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_2_impl_out,
                 X => Delay1No140_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast);

Delay7No82_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast <= Delay7No82_out;
SharedReg439_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg439_out;
SharedReg258_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg258_out;
SharedReg461_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg461_out;
SharedReg39_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg9_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg473_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg473_out;
SharedReg449_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg449_out;
SharedReg415_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg415_out;
SharedReg260_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg475_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg475_out;
SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg6_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
   MUX_Product102_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No82_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg439_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg475_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg258_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg461_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg473_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg449_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg415_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product102_2_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_0_out,
                 Y => Delay1No140_out);

SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg31_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg393_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg393_out;
   MUX_Product102_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg572_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg569_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg393_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg573_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg568_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product102_2_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product431_0_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product431_0_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product431_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product431_0_impl_out,
                 X => Delay1No142_out_to_Product431_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product431_0_impl_parent_implementedSystem_port_1_cast);

SharedReg221_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg24_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg9_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg190_out;
SharedReg445_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg445_out;
SharedReg466_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg466_out;
SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg458_out;
SharedReg459_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg459_out;
SharedReg351_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg351_out;
SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg458_out;
SharedReg365_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg190_out;
   MUX_Product431_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg351_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg190_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg445_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg466_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg458_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg459_out_to_MUX_Product431_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product431_0_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_0_impl_0_out,
                 Y => Delay1No142_out);

SharedReg567_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg32_out;
SharedReg4_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg571_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg17_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg364_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg364_out;
SharedReg23_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg23_out;
SharedReg573_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg573_out;
   MUX_Product431_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg364_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg23_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg573_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg32_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product431_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product431_0_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_0_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Product431_1_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Product431_1_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Product431_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product431_1_impl_out,
                 X => Delay1No144_out_to_Product431_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Product431_1_impl_parent_implementedSystem_port_1_cast);

SharedReg373_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg282_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg168_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg195_out;
SharedReg24_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg9_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg195_out;
SharedReg461_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg461_out;
SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg473_out;
SharedReg451_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg451_out;
SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg473_out;
SharedReg28_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg28_out;
   MUX_Product431_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg451_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg473_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg195_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg461_out_to_MUX_Product431_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product431_1_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_1_impl_0_out,
                 Y => Delay1No144_out);

SharedReg394_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg23_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg573_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg32_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg32_out;
SharedReg570_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
SharedReg372_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Product431_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg32_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg573_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product431_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product431_1_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_1_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product481_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product481_2_impl_out,
                 X => Delay1No146_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast);

SharedReg177_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg482_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg482_out;
SharedReg28_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg319_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg291_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg174_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg174_out;
SharedReg201_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg201_out;
SharedReg24_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg9_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg236_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg236_out;
SharedReg507_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg507_out;
SharedReg562_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg562_out;
   MUX_Product481_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg482_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg236_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg507_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg28_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg174_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg201_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product481_2_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_2_impl_0_out,
                 Y => Delay1No146_out);

SharedReg570_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg318_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg379_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg23_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg573_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg31_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
   MUX_Product481_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg573_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product481_2_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_2_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product491_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product491_0_impl_out,
                 X => Delay1No148_out_to_Product491_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product491_0_impl_parent_implementedSystem_port_1_cast);

SharedReg445_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg445_out;
SharedReg1_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg221_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg221_out;
SharedReg458_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg458_out;
SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg459_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg459_out;
SharedReg466_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg466_out;
SharedReg28_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg406_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg365_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg252_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg252_out;
   MUX_Product491_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg445_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg252_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg221_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg458_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg459_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg466_out_to_MUX_Product491_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product491_0_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_0_impl_0_out,
                 Y => Delay1No148_out);

SharedReg567_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg405_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg405_out;
SharedReg352_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg352_out;
SharedReg36_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg36_out;
SharedReg573_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg573_out;
   MUX_Product491_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg405_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg36_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg573_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg559_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product491_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product491_0_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_0_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product491_1_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product491_1_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product491_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product491_1_impl_out,
                 X => Delay1No150_out_to_Product491_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product491_1_impl_parent_implementedSystem_port_1_cast);

SharedReg281_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg281_out;
SharedReg282_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg229_out;
SharedReg258_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg258_out;
SharedReg1_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg229_out;
SharedReg473_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg473_out;
SharedReg562_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg171_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg171_out;
SharedReg439_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg439_out;
SharedReg280_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg280_out;
   MUX_Product491_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg281_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg171_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg439_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg280_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg258_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg229_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg473_out_to_MUX_Product491_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product491_1_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_1_impl_0_out,
                 Y => Delay1No150_out);

SharedReg373_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg36_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg573_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg570_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
SharedReg393_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg393_out;
   MUX_Product491_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg393_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg573_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg559_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product491_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product491_1_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_1_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product512_0_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product512_0_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product512_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_0_impl_out,
                 X => Delay1No152_out_to_Product512_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product512_0_impl_parent_implementedSystem_port_1_cast);

SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg458_out;
SharedReg38_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg9_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg458_out;
SharedReg252_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg252_out;
SharedReg466_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg466_out;
SharedReg433_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg433_out;
SharedReg163_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg163_out;
SharedReg498_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg498_out;
SharedReg363_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg363_out;
SharedReg364_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg364_out;
SharedReg499_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg499_out;
SharedReg435_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg435_out;
   MUX_Product512_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg363_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg364_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg499_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg435_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg458_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg252_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg466_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg433_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg163_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg498_out_to_MUX_Product512_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_0_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_0_impl_0_out,
                 Y => Delay1No152_out);

SharedReg567_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg25_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg570_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg351_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg351_out;
SharedReg406_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg565_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg565_out;
SharedReg566_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg566_out;
   MUX_Product512_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg351_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg565_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg566_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg568_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product512_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_0_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_0_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product512_1_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product512_1_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product512_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_1_impl_out,
                 X => Delay1No154_out_to_Product512_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product512_1_impl_parent_implementedSystem_port_1_cast);

SharedReg394_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg474_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg474_out;
SharedReg440_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg440_out;
SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg449_out;
SharedReg38_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg38_out;
SharedReg9_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg461_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg461_out;
SharedReg258_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg258_out;
SharedReg439_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg439_out;
SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg415_out;
SharedReg198_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg198_out;
SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg415_out;
SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg449_out;
   MUX_Product512_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg474_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg198_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg415_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg440_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg449_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg38_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg461_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg258_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg439_out_to_MUX_Product512_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_1_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_1_impl_0_out,
                 Y => Delay1No154_out);

SharedReg373_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg565_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg565_out;
SharedReg566_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg25_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg570_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg564_out;
   MUX_Product512_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg565_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg564_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg566_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg568_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Product512_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_1_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_1_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product512_2_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product512_2_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product512_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_2_impl_out,
                 X => Delay1No156_out_to_Product512_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product512_2_impl_parent_implementedSystem_port_1_cast);

SharedReg203_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg507_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg507_out;
SharedReg289_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg289_out;
SharedReg290_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg290_out;
SharedReg291_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg236_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg236_out;
SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg1_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg2_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg263_out;
SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg422_out;
   MUX_Product512_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg507_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg422_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg289_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg290_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg291_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg236_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product512_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_2_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_2_impl_0_out,
                 Y => Delay1No156_out);

SharedReg570_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg378_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg378_out;
SharedReg319_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg36_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg573_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg560_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg3_out;
   MUX_Product512_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg3_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg378_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg573_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product512_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_2_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_2_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product512_3_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product512_3_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product512_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_3_impl_out,
                 X => Delay1No158_out_to_Product512_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product512_3_impl_parent_implementedSystem_port_1_cast);

SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg265_out;
SharedReg516_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg516_out;
SharedReg562_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg562_out;
SharedReg182_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg488_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg488_out;
SharedReg28_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg327_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg335_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg179_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg179_out;
SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg265_out;
SharedReg24_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg2_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg558_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product512_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg516_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg562_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg182_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg488_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg179_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg265_out_to_MUX_Product512_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_3_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_3_impl_0_out,
                 Y => Delay1No158_out);

SharedReg560_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg562_out;
SharedReg570_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg326_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg386_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg23_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg573_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg20_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg559_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg559_out;
   MUX_Product512_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg559_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg562_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg573_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product512_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_3_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_3_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product512_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_4_impl_out,
                 X => Delay1No160_out_to_Product512_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product512_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg492_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg492_out;
SharedReg184_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg184_out;
SharedReg524_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg524_out;
SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg540_out;
SharedReg493_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg493_out;
SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg540_out;
SharedReg28_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg344_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg344_out;
SharedReg525_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg525_out;
SharedReg155_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg155_out;
SharedReg267_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg267_out;
SharedReg38_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg38_out;
SharedReg2_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
   MUX_Product512_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg492_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg155_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg267_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg38_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg184_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg524_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg493_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg540_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg344_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg525_out_to_MUX_Product512_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_4_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_4_impl_0_out,
                 Y => Delay1No160_out);

SharedReg558_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg343_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg343_out;
SharedReg401_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg401_out;
SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg565_out;
SharedReg573_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg556_out;
SharedReg25_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Product512_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg573_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg556_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg563_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg343_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg401_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg565_out_to_MUX_Product512_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product512_4_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_4_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product611_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_0_impl_out,
                 X => Delay1No162_out_to_Product611_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product611_0_impl_parent_implementedSystem_port_1_cast);

SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg466_out;
SharedReg39_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg9_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg466_out;
SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg445_out;
SharedReg498_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg498_out;
SharedReg253_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg253_out;
SharedReg194_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg194_out;
SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg433_out;
SharedReg458_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg458_out;
SharedReg352_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg352_out;
SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg433_out;
SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg445_out;
   MUX_Product611_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg458_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg466_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg445_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg498_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg253_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg194_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg433_out_to_MUX_Product611_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_0_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_0_impl_0_out,
                 Y => Delay1No162_out);

SharedReg567_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg31_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg564_out;
SharedReg406_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg572_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg573_out;
   MUX_Product611_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg564_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg572_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg573_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg31_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg568_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg569_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product611_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_0_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_0_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product611_2_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product611_2_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product611_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_2_impl_out,
                 X => Delay1No164_out_to_Product611_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product611_2_impl_parent_implementedSystem_port_1_cast);

SharedReg510_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg510_out;
SharedReg422_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg422_out;
SharedReg263_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg379_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg483_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg483_out;
SharedReg508_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg508_out;
SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg453_out;
SharedReg38_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg38_out;
SharedReg9_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg482_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg482_out;
SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg453_out;
SharedReg98_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg98_out;
SharedReg264_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg264_out;
   MUX_Product611_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg510_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg422_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg482_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg98_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg264_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg263_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg483_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg508_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg453_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg38_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product611_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_2_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_2_impl_0_out,
                 Y => Delay1No164_out);

SharedReg570_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg319_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg565_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg566_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg556_out;
SharedReg25_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg569_out;
   MUX_Product611_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg568_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg561_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg569_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg564_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg566_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg556_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg558_out_to_MUX_Product611_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_2_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_2_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product611_3_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product611_3_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product611_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_3_impl_out,
                 X => Delay1No166_out_to_Product611_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product611_3_impl_parent_implementedSystem_port_1_cast);

SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg488_out;
SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg532_out;
SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg532_out;
SharedReg211_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg211_out;
SharedReg516_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg516_out;
SharedReg333_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg333_out;
SharedReg334_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg334_out;
SharedReg335_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg243_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg243_out;
SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg488_out;
SharedReg1_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg9_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg488_out;
   MUX_Product611_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg532_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg211_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg516_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg333_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg334_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg243_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg488_out_to_MUX_Product611_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_3_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_3_impl_0_out,
                 Y => Delay1No166_out);

SharedReg560_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg3_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg570_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg385_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg385_out;
SharedReg327_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg36_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg36_out;
SharedReg573_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg25_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg558_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
   MUX_Product611_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg3_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg385_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg36_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg573_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product611_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_3_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_3_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product611_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product611_4_impl_out,
                 X => Delay1No168_out_to_Product611_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product611_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg524_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg524_out;
SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg216_out;
SharedReg540_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg540_out;
SharedReg248_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg248_out;
SharedReg131_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg131_out;
SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg555_out;
SharedReg307_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg307_out;
SharedReg308_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg555_out;
SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg216_out;
SharedReg492_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg492_out;
SharedReg39_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg39_out;
SharedReg9_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg9_out;
   MUX_Product611_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg524_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg492_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg39_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg216_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg540_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg248_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg131_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg307_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg555_out_to_MUX_Product611_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_4_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_4_impl_0_out,
                 Y => Delay1No168_out);

SharedReg558_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg400_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg400_out;
SharedReg344_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg344_out;
SharedReg572_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg573_out;
SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg556_out;
SharedReg25_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Product611_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg573_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg556_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg560_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg569_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg563_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg400_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg344_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg572_out_to_MUX_Product611_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product611_4_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product611_4_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product811_3_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product811_3_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product811_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product811_3_impl_out,
                 X => Delay1No170_out_to_Product811_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product811_3_impl_parent_implementedSystem_port_1_cast);

SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg516_out;
SharedReg427_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg427_out;
SharedReg245_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg534_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg534_out;
SharedReg532_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg532_out;
SharedReg265_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg265_out;
SharedReg386_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg517_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg517_out;
SharedReg533_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg533_out;
SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg516_out;
SharedReg38_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg38_out;
SharedReg9_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg558_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg516_out;
   MUX_Product811_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg427_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg38_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg245_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg534_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg532_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg265_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg517_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg533_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg516_out_to_MUX_Product811_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product811_3_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_3_impl_0_out,
                 Y => Delay1No170_out);

SharedReg560_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg561_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg569_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg570_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg563_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg564_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg564_out;
SharedReg327_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg327_out;
SharedReg565_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg566_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg556_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg556_out;
SharedReg31_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg558_out;
SharedReg568_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg568_out;
   MUX_Product811_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg556_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg558_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg568_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg564_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg327_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg566_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Product811_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product811_3_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_3_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product811_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product811_4_impl_out,
                 X => Delay1No172_out_to_Product811_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product811_4_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg40_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg158_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg158_out;
SharedReg269_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg269_out;
SharedReg524_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg524_out;
SharedReg540_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg540_out;
SharedReg267_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg267_out;
SharedReg555_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg555_out;
SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg541_out;
SharedReg247_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg247_out;
SharedReg401_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg401_out;
SharedReg558_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg558_out;
   MUX_Product811_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg401_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg558_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg158_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg269_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg524_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg540_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg267_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg555_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg541_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg247_out_to_MUX_Product811_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product811_4_impl_0_LUT_out,
                 oMux => MUX_Product811_4_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_4_impl_0_out,
                 Y => Delay1No172_out);

SharedReg31_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg344_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg561_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg561_out;
SharedReg560_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg560_out;
SharedReg558_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg558_out;
SharedReg570_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg569_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg569_out;
SharedReg567_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg568_out;
SharedReg564_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg566_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg566_out;
SharedReg556_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg556_out;
   MUX_Product811_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg566_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg561_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg560_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg558_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg569_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg567_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg568_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Product811_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product811_4_impl_1_LUT_out,
                 oMux => MUX_Product811_4_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product811_4_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Subtract12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_0_impl_out,
                 X => Delay1No174_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast);

Delay72No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast <= Delay72No_out;
SharedReg235_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg235_out;
SharedReg42_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg42_out;
SharedReg193_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg193_out;
SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg44_out;
SharedReg74_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg74_out;
SharedReg165_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg165_out;
SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg44_out;
SharedReg166_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg166_out;
SharedReg113_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg113_out;
SharedReg227_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg227_out;
SharedReg164_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg164_out;
SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg228_out;
SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg224_out;
   MUX_Subtract12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay72No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg235_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg227_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg164_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg42_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg193_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg74_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg165_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg44_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg166_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg113_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_0_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_0_out,
                 Y => Delay1No174_out);

SharedReg355_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg355_out;
SharedReg283_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg283_out;
SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg405_out;
SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg271_out;
SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg271_out;
SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg405_out;
SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg271_out;
SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg365_out;
SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg365_out;
SharedReg272_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg272_out;
SharedReg369_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg369_out;
   MUX_Subtract12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg355_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg283_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg272_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg369_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg405_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg271_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg365_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_0_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Subtract12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_1_impl_out,
                 X => Delay1No176_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg172_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg172_out;
SharedReg87_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg87_out;
SharedReg232_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg232_out;
Delay72No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast <= Delay72No1_out;
SharedReg207_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg207_out;
SharedReg434_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg434_out;
SharedReg170_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg170_out;
SharedReg436_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg436_out;
SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg51_out;
SharedReg140_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg140_out;
SharedReg52_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg52_out;
SharedReg141_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg141_out;
SharedReg82_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg82_out;
SharedReg200_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg200_out;
   MUX_Subtract12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg172_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg52_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg141_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg82_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg200_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg232_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay72No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg207_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg434_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg170_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg436_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg51_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg140_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_1_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_0_out,
                 Y => Delay1No176_out);

SharedReg282_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg320_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg320_out;
SharedReg377_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg293_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg293_out;
SharedReg292_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg292_out;
SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg393_out;
SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg280_out;
SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg280_out;
SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg393_out;
SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg280_out;
SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg374_out;
SharedReg376_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg376_out;
   MUX_Subtract12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg320_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg374_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg376_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg377_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg293_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg292_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg393_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg280_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_1_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Subtract12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_2_impl_out,
                 X => Delay1No178_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast);

Delay13No12_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast <= Delay13No12_out;
SharedReg127_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg127_out;
Delay29No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast <= Delay29No2_out;
SharedReg178_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg92_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg92_out;
SharedReg204_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg204_out;
Delay72No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast <= Delay72No2_out;
Delay32No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast <= Delay32No3_out;
SharedReg416_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg416_out;
SharedReg143_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg143_out;
SharedReg418_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg418_out;
SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg58_out;
SharedReg122_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg122_out;
SharedReg59_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg59_out;
   MUX_Subtract12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay13No12_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg418_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg58_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg122_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg59_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay29No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg92_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg204_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay72No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay32No3_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg416_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg143_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_2_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_0_out,
                 Y => Delay1No178_out);

SharedReg320_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg320_out;
SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg383_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg383_out;
SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg291_out;
SharedReg335_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg335_out;
SharedReg384_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg384_out;
SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg303_out;
SharedReg302_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg302_out;
SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg300_out;
SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg318_out;
SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg318_out;
SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg300_out;
SharedReg289_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg289_out;
SharedReg380_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg380_out;
   MUX_Subtract12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg320_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg289_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg380_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg383_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg291_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg335_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg384_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg303_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg302_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg300_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg318_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract12_2_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Subtract12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_4_impl_out,
                 X => Delay1No180_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg159_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg159_out;
SharedReg69_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg105_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg160_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg160_out;
Delay9No24_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast <= Delay9No24_out;
SharedReg186_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg186_out;
SharedReg132_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg132_out;
Delay32No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast <= Delay32No4_out;
Delay72No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast <= Delay72No4_out;
   MUX_Subtract12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg159_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg105_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg160_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay9No24_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg186_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay32No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay72No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Subtract12_4_impl_0_LUT_out,
                 oMux => MUX_Subtract12_4_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_4_impl_0_out,
                 Y => Delay1No180_out);

SharedReg307_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg307_out;
SharedReg343_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg343_out;
SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg310_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg310_out;
SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg345_out;
SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg400_out;
SharedReg309_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg309_out;
SharedReg404_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg404_out;
   MUX_Subtract12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg343_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg310_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg345_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg309_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg404_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Subtract12_4_impl_1_LUT_out,
                 oMux => MUX_Subtract12_4_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_4_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Subtract1_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract1_3_impl_out,
                 X => Delay1No182_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast);

SharedReg63_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg64_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
Delay13No13_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast <= Delay13No13_out;
SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg183_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg183_out;
SharedReg152_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg152_out;
SharedReg189_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg189_out;
SharedReg212_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg212_out;
Delay72No3_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast <= Delay72No3_out;
SharedReg188_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg188_out;
SharedReg99_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg99_out;
SharedReg150_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg150_out;
SharedReg102_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg102_out;
   MUX_Subtract1_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg188_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg99_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg150_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg102_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg64_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay13No13_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg183_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg152_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg189_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg212_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay72No3_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract1_3_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_3_impl_0_out,
                 Y => Delay1No182_out);

SharedReg385_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg385_out;
SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg307_out;
SharedReg328_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg328_out;
SharedReg335_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg335_out;
SharedReg345_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg345_out;
SharedReg330_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg330_out;
SharedReg301_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg301_out;
SharedReg346_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg346_out;
SharedReg392_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg392_out;
SharedReg390_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg390_out;
SharedReg348_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg348_out;
SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg307_out;
SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg333_out;
SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg333_out;
   MUX_Subtract1_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg385_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg348_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg307_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg333_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg328_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg335_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg345_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg330_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg301_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg346_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg392_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg390_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract1_3_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_3_impl_1_out,
                 Y => Delay1No183_out);
   Constant1_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

Delay1No184_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Divide_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_0_impl_out,
                 X => Delay1No184_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast);

SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg552_out;
SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg552_out;
SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg552_out;
SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg552_out;
SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg552_out;
   MUX_Divide_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg552_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Divide_0_impl_0_LUT_out,
                 oMux => MUX_Divide_0_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_0_out,
                 Y => Delay1No184_out);

SharedReg405_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg405_out;
SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg318_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg326_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg326_out;
SharedReg400_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg400_out;
   MUX_Divide_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg405_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg318_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg326_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg400_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Divide_0_impl_1_LUT_out,
                 oMux => MUX_Divide_0_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product45_4_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product45_4_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product45_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product45_4_impl_out,
                 X => Delay1No186_out_to_Product45_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product45_4_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg31_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg247_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg247_out;
SharedReg542_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg542_out;
SharedReg267_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg267_out;
   MUX_Product45_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg247_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg542_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Product45_4_impl_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Product45_4_impl_0_LUT_out,
                 oMux => MUX_Product45_4_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product45_4_impl_0_out,
                 Y => Delay1No186_out);

SharedReg14_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg400_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg570_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg573_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg573_out;
SharedReg560_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg560_out;
   MUX_Product45_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg570_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg573_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg560_out_to_MUX_Product45_4_impl_1_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Product45_4_impl_1_LUT_out,
                 oMux => MUX_Product45_4_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product45_4_impl_1_out,
                 Y => Delay1No187_out);
   Constant_0_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);

   Delay156No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => Delay156No_out);

   Delay156No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => Delay156No1_out);

   Delay156No4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => Delay156No4_out);

   Delay145No3_instance: Delay_34_DelayLength_133_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=133 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => Delay145No3_out);

   Delay151No_instance: Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=139 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay151No_out);

   Delay151No1_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => Delay151No1_out);

   Delay151No2_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => Delay151No2_out);

   Delay151No3_instance: Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=139 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => Delay151No3_out);

   Delay151No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => Delay151No4_out);

   Delay154No7_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay154No7_out);

   Delay154No8_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => Delay154No8_out);

   Delay156No5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay156No5_out);

   Delay156No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => Delay156No6_out);

   Delay156No9_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => Delay156No9_out);

   Delay22No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay22No_out);

   Delay22No1_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => Delay22No1_out);

   Delay22No4_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => Delay22No4_out);

   Delay13No5_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay13No5_out);

   Delay13No6_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => Delay13No6_out);

   Delay11No5_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => Delay11No5_out);

   Delay11No7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay11No7_out);

   Delay11No8_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay11No8_out);

   Delay9No24_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => Delay9No24_out);

   Delay16No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => Delay16No_out);

   Delay16No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => Delay16No1_out);

   Delay16No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => Delay16No2_out);

   Delay16No3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => Delay16No3_out);

   Delay16No4_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => Delay16No4_out);

   Delay13No12_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => Delay13No12_out);

   Delay13No13_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => Delay13No13_out);

   Delay32No3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => Delay32No3_out);

   Delay32No4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => Delay32No4_out);

   Delay22No5_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => Delay22No5_out);

   Delay22No6_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => Delay22No6_out);

   Delay22No9_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => Delay22No9_out);

   Delay18No11_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => Delay18No11_out);

   Delay29No2_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => Delay29No2_out);

   Delay7No82_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => Delay7No82_out);

   Delay7No83_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => Delay7No83_out);

   Delay2No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => Delay2No120_out);

   Delay2No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => Delay2No121_out);

   Delay2No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => Delay2No122_out);

   Delay2No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => Delay2No123_out);

   Delay2No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => Delay2No124_out);

   Delay12No39_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => Delay12No39_out);

   Delay82No_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => Delay82No_out);

   Delay82No1_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => Delay82No1_out);

   Delay82No4_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => Delay82No4_out);

   Delay88No_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => Delay88No_out);

   Delay88No1_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => Delay88No1_out);

   Delay88No2_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => Delay88No2_out);

   Delay88No3_instance: Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=80 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => Delay88No3_out);

   Delay88No4_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => Delay88No4_out);

   Delay130No5_instance: Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=122 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => Delay130No5_out);

   Delay130No6_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => Delay130No6_out);

   Delay130No7_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => Delay130No7_out);

   Delay130No8_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => Delay130No8_out);

   Delay130No9_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => Delay130No9_out);

   Delay73No_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => Delay73No_out);

   Delay73No3_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => Delay73No3_out);

   Delay72No_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => Delay72No_out);

   Delay72No1_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => Delay72No1_out);

   Delay72No2_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => Delay72No2_out);

   Delay72No3_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => Delay72No3_out);

   Delay72No4_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => Delay72No4_out);

   Delay42No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => Delay42No_out);

   Delay42No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => Delay42No1_out);

   Delay42No2_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => Delay42No2_out);

   Delay41No2_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => Delay41No2_out);

   Delay45No_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => Delay45No_out);

   Delay45No1_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => Delay45No1_out);

   Delay45No2_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => Delay45No2_out);

   Delay45No3_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => Delay45No3_out);

   Delay45No4_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay45No4_out);

   Delay34No4_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => Delay34No4_out);

   Delay116No1_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => Delay116No1_out);

   Delay116No2_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => Delay116No2_out);

   Delay116No3_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => Delay116No3_out);

   Delay116No4_instance: Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=115 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => Delay116No4_out);

   Delay118No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => Delay118No_out);

   Delay118No1_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => Delay118No1_out);

   Delay118No2_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => Delay118No2_out);

   Delay118No3_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => Delay118No3_out);

   Delay118No4_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => Delay118No4_out);

   MUX_Inv_11_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_11_0_0_LUT_out);

   MUX_Inv_12_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_12_0_0_LUT_out);

   MUX_Inv_13_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_13_0_0_LUT_out);

   MUX_Inv_21_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_21_0_0_LUT_out);

   MUX_Inv_22_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_22_0_0_LUT_out);

   MUX_Inv_23_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_23_0_0_LUT_out);

   MUX_Inv_31_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_31_0_0_LUT_out);

   MUX_Inv_32_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_32_0_0_LUT_out);

   MUX_Inv_33_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_33_0_0_LUT_out);

   MUX_Inv_41_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_41_0_0_LUT_out);

   MUX_Inv_42_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_42_0_0_LUT_out);

   MUX_Inv_43_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Inv_43_0_0_LUT_out);

   MUX_Add31_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add31_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Add31_4_impl_0_LUT_out);

   MUX_Add31_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add31_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Add31_4_impl_1_LUT_out);

   MUX_Product811_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product811_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product811_4_impl_0_LUT_out);

   MUX_Product811_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product811_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product811_4_impl_1_LUT_out);

   MUX_Subtract12_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract12_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Subtract12_4_impl_0_LUT_out);

   MUX_Subtract12_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract12_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Subtract12_4_impl_1_LUT_out);

   MUX_Divide_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Divide_0_impl_0_LUT_out);

   MUX_Divide_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Divide_0_impl_1_LUT_out);

   MUX_Product45_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product45_4_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product45_4_impl_0_LUT_out);

   MUX_Product45_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product45_4_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product45_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_0_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_0_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_0_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_0_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_0_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_1_impl_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_2_impl_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_3_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_4_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_0_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_1_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_2_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_3_impl_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_4_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_3_impl_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_4_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_0_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_1_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_2_impl_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_3_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_4_impl_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_0_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_1_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_2_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_3_impl_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_4_impl_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_0_impl_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_1_impl_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_2_impl_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_3_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_4_impl_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_0_impl_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_1_impl_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_2_impl_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_3_impl_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_4_impl_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_0_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_1_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_2_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_3_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_4_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_0_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_1_impl_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_2_impl_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_3_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_4_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_0_impl_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=117 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_1_impl_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=117 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_2_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=137 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_3_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_119_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=119 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_4_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=117 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_2_impl_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=115 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_3_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_120_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=120 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_3_impl_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_136_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=136 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_4_impl_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=115 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_1_impl_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=117 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_0_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=115 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_1_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_2_impl_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_3_impl_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_2_impl_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=124 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_4_impl_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_0_impl_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add31_4_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_139_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=139 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_2_impl_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_3_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_4_impl_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_1_impl_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_2_impl_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product431_0_impl_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product431_1_impl_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product481_2_impl_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product491_0_impl_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product491_1_impl_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_0_impl_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_1_impl_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_2_impl_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_3_impl_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_4_impl_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_0_impl_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_2_impl_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_3_impl_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product611_4_impl_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product811_3_impl_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product811_4_impl_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_0_impl_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_1_impl_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_2_impl_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_4_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract1_3_impl_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_165_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=165 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_0_impl_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product45_4_impl_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);
end architecture;

